PK   Pn5[I幯�  �;     cirkitFile.json�Z[s�:�+�j��qQ����n��LR����8�AĜ����lj��J��U��rbԭ�[�SwK�f�Ef�0/��Ee�g�vg�Zѫ8nE3{�d�*_>b��o���S��J'�7�<�Y�.�E��&�tV���s!�*��Ⱦy����E��!H�����D��«�eKb?ͮ��!��2Q��)�;�uwa�=Xw�=�u��0YA넂Lc�M�d��i�a�S�mX|.4<��&�(��F>��0a&Fu��C�y�:��2�i1�!�k��n3z��y���.
������| 
�Q� �AaFP\#(��J`�k�8�."���E��C`��1ᆾnL9���1C`|��S��x|����B.E���g�zS���:����ҥ������L�B��� G!FP�f�5��A�FP��"��b3��f���_d��� G�8O�S��,MNp��9R�!�?���a�D?�wf�&�,��T�2Z�̑�T;�G�i$[<� '��[FC���a ���ɧ\��PL|z:Я���E�OdQ���7>>i� ��u��N�@��`�j��"�%Y[[��y�m�K"hٍN?���9dA������������}`� ؟���2z�
:����ե�;���6�%0a��{Z@�\yC��/ȉJ�tA�V���2�_�B��D:g(�R'�)����ۤǦҔt��S_}���ιu��Zk�:b��h������i 1��Ù�+W�	D� >����F���~����@���NgD=��;�iz��9'1�alwr�@Ͽ`��p{b�;fWzs���L5�ϙm���g�g���H#"�"ڈ蹈5"�#�H�媐"Z�ZU۪8_�IY��߰���GQ	��V7��VU"u�҇�y�T�kF����s)����Mq@����U�c�E��D��G�9>����,�ƞ`��o�M3[�Jd�hR���y�(����m5vR��l��ȸ?wg�#�������9�sݮs���mnp'��\���\��^���E^m�g��N ��k⵶2�]�(�|`���s�)G���5��1sZ��5O�1B���5��g@��0.%rR�xA0 GuJ���L�Yp༯�gjr$�C����厍�tN�R�!���f��f��,�"ɞK2���Z:�_D��W?}s0
�vY�։�~����.�U��M,�R*a)�oI��Rٶ�߻����U��j�lD��EX�
Y��p����ŏ�2��.b5_s�&�u�?�"2�c���k���5���"��;""��sB)����J'��I�Ȅ5M=�״�yE�Z@�ޡ���cތ� �{M��nh߃�(	���k0h-��j�6j8#8hts�]Zk�"�*�J���m��gֿ�~�DY���4��-��Bl6��?�\D�-̣�s�gU���,��q�0�uRZIe)"���ZI+JJ��ɰ��煕��F��C=V[��)qn��r��3�o�TI��h�mS;ܣ�f�:�r���̎�d{{��}~O��}k�Y���s�����M�T��{�n>��g|�]���OG�g�՚�������y����^Ǌ�d/j+�|$���\��a���1�N���霩��U2���ľZk��G*�����E('�+�*��:���	��xZ�����.]�iZԁ�ʷZ�9i�0���G,P��nzM�j��0э���Z&�k�HU_����ӎ�N���T�k�������_���]����ma������n�-T �Zv��]����d�BM+�k�B�>�tM�}2��6OT�պ�z[,�����{-x��B�[o��:ɵ�R�yW�k�Y���b�Z�>��
��jk�-�k=�^ؿ}O����$�9*"�T$F����⡤"�T|��O���8�kQ�K2ϿB��k�Z�Tܿf���`T4�Ej6,^Gƶ�w���Nk�f؟B�wZ�W����[�>-���.���C��֟h��{����e�$��9bsüfFyͯ�u�	��;�¢I1��ꍋ�B�9�D��Zݡ� �ϴ�u���DZO<!6��tb��Elz��OUw.x2����D��r�gZ{r��W��w�Q�"���h�����G_D����s%7�~Υ�&�_2�>�2,�m����PK   Pn5[����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   Pn5[԰�B� .4 /   images/44d6884f-a329-4b4e-966d-57539d09419f.png�|eXT]�� H;�"]�%a���
�ҥ�HH�t �H�� �9(HC��������x�|��}�]k�u�y��ڋ��SMe��L!���c�t	![�$Zn��T �.��y@ ��$��Hj���S񙧮����wk����������Wkw۴��L�-���z��W��zx�����Ka#�[H�R���(��[��H߱TG�c0�U[��//G��<�P��@�F]��ӧt$��I���_�u�nJJ��1I�-U������U�=����HXa�@fq'��B���h���FQn���7��U���	�2.��ӪL�`��UO3��;��yz��]&���a�^?X\s���<��	_�ݱ����˫��B����Y�3�T>��>�R(� ���hі$�_Zf�c�#��*ڷ���"?b{E� [~P���+�č"�����%E�~��+���w��jCЕw�Hͭ5kr<�xL��~�>9m:!����� �K�8'y��@;����&�,Ǝ'Ւ
_P���s��g���1w0�kə���W@��^T�'�P��Y�}�qoұٸ���<f@<��
!����'88o���v���U��;�fS�"�gRRRВ��!S��+d	�D��T�7
��,�a���&h�ͽ�@�x�柷�eϪ,���H !R���0�sY��V��rUB�{3�N���X����RRR���a��h��󪝉��;�!~�k�����]���Ľ5�A�V�3V��8}p`c2x^F�Ż0	t�>�x%@n&��gC����RE��>za�E+�	D`L�|��ɳ<i����ynAA-
�O����WE|Q�*H2��@|��S�5a4���q]]]��7���ITf�����D�4��%�6L�&,���|�z�������17�O��;��}}}�0���X�n0Z�1[ѹ`0�<fw��KFFF�I���'q���ӡ$�7���,l��q�	���G�����`�MpY��C7�<}Z�9HEV:A�i�DOS��<�"�6-��3c���HZ|�qMX�������X�׆�\GFF�1�X���(�Λ��k?00�� d{h��B\og�aƟ��m�Wf4:����Y��ڟ��u��]n��c�%e��Տ7��~��A�\p;5@����+q�;Uxb�̫�ОR�sp�r'ՍgI�Q�)���&����i�.�P'dR.@H�T�w@��qt��Ѩ �[�6�3\�A�tL����\��>R�IS�'�=�)J��	j���/�B�8lR�n�Fs4��!k������鳋og�18qQ����_����̺�� ��xά�s��>�U=Űl�f����57g9��H�V>��д�^�>Um�ի"�R�>�����8�\������FT#UT����k@�����ۃ��ۏ'g�!7T$�Wq�c|��� ��C鹬;u��?�"��fj m�*�.\��411���姨c>�B-�{����3��+�k��.]�i���?����.�����QX���v�[Aef�v��>'$�| �����\%���Ezz�>q��|($���' W>v1�>-4�p�1g�I���􇛣&����g?�\���<�"����v2�.@��ذ�+(|��Bz�><��qc6399���谘r������p�H�L/ZW�Dp��R����'�}����G�c~#��<�_ð��;��þ5oǿ�+�,��SـKt0�,#�W�2����4HA��7�c9��e����<͜z
ȭ#�����v�����J*���\z�gl�2߳y���t�r�wC���iwjj�v�t§�Wnى�Tҩ�D���s�1~l����[����a���x.�g�/ڕ�<�u�\�%�����0�I�9�����g�|��"�o���glPyQ�� �S������:����z�{u|�M�(���\���-���@�J >wvt����[�lk[�W��!��Z	�I�� �7o�XH�Wi���lL����̪n�iMx���2EԪ[��k%i^��9?����@u�_��)�y�k�0�C��Z���l�z!t5ߊK|�w6+�IM	A?&3�Z
�<�ת;���Yo����4�|���ſ�|��y�v֕-�FMOO�n��̶���P����^cJ����Z�1�P:J.Sf+�$kԭbX����o�u�̎� *��If�d������с�!tN*FF�su�$�@�9a�t�zΦ�[�����e���0���+��^�=My���`��@��+�����ΌR-ث�2ԊXS���.�� �N��f�Q����߼�c���w�_��_���g#�@��3Tz�Js����R�����{�T���������B�W�8��������x咈��-.�z#-��sg
�������O�L�-�B��ޣ�L͢;C��Z�R��N�� st2XU7�o�𲅽!�Q��=����uI�5�.y����m�{�l�t��fc�^������i"`cR��QP2:�F�W(��;`�u��O�0c;����#���L�~ ��:E�q��s�U�����,�~ P�񳭃�g��Z��FcAĴB2`m���Y;����L���E�^�Ϭ��2JJ���t�c�k�u��	��hW`�ѿ�Mn��@��6��2��
_nҐ �|]��O�������r^�:�O��h\ҿ��� 2��
j����>��K����9��K"ք��)�#;��}5��Jf���@p�d�������>�l�A�~��ׇ��jQ1����}{�2h�+V����UulllJ�2��P~gd��<�y���9���/(8V�_Z�#���Tnt�//��4K���\%Ua��9��x�� l���<��� D��ځ�y��H��Dv�?��6��ޤ�~
%=�\;���%9:�U)�g���g�^�/i��E�lp��������#/�̏c���#��ˍ5�$T�v����W�K@J����9��s.�H�qΠ�v<���uq��V�0�$�0���h� 5r�pCL�����_�w��<選
q��0���iY	y����N�Z��]��_��vƖU�ޭ�p�@�u��[�a�BF߆�������o���J��� 8��/�|oz&�#5��T����_���@��f?�����\�,��y�$�3`�s� j�ѻ��D�� A�r/��݀���`o�?��_�V�[@�HBI�
�U��t�>'Riu������ڙ�C���P���9�'�l![6)�L��!Me����(cP�ı�D&��s�����;	�A{6u8���p0v�ʀRY�K���w�F)��v��>�9�Zpy�s�w��{���L��_A�����8�u��� ذ`w�]P**泝y�s0��Z���(�3(U뙞���"�y��������S�?�i����ά����\��T�+���,����g��i�c���-bG��_�����?���%�5��+���)%m�����B�l�!@��Fs�&ƓTJ�c�2���(��?�'l��<���wZ|ýzn
(�M�)P.�Rgp��r[Y�s:a�kXBA���;H%*�f`�l�·���NE�5ܠ�᷺��'�7�M4�r���:�A˟���~���oj��u���퇊���.� aʾ\.���.1!�`�L�ڦFW��q�)Uֳ������k��e?��&�=Fn�2�I���t����3� �.ò����9Y �V_�� Oa�]+x\�#.�~t4�Tn-�ړw��q5������?3V=�J�����	�+������E�������ݑ��nk*nX.�ݎV*Պ���H(���y��w�%������MI�H��?f�a6Y�u�E�6Y���\��]l����s����3��
K�H���`3��h��[�3L
����4��Ɍ�|�^��2WXDD����Q�cEE�8�Kx�3\jZ�Ԫ���|�Z3��1����\��s�A��;N�p��ҼK��Z_�{YQ��!�˺�p_7�J ^���R�[�%ojDu�J-�1G�uT��\�s��u��&q��p��/ʱ�:����n:ZZTĥ�p��a� �C#5o�"،��=Ι�S�%!�q�o[b��,C�977�ò=B���;�4Y��رy�X�b#�So�[2-$k�EyOo_ ���Rv �T�^*��S�g��ؤ8?��r��돶�33Y��3�ǟQA��G˴��R�Đ0LAI�Z4�|��2�:��d��̃��
�$H�xܴ����Sc���3��"�R)�L�YM��G��\ʵK!,�4�Bl�vK��������~`�79�X�*�;�W� ��H2�S�����dm����沋Ns�ūh?hd#�(��/,,�j���C���aW��>���z���S����s�{��R#t;��y��c��!�v�CgX�<�,���]��_����S�%��j�~��)/S�_�>�@��G���Z���-5��ɕ�	�}K�zm��z3d�����aΛI:��u||�z'�+�4��.#�툴��=W�e���C�u��呛�.{;���7�E3���H%g�M����Qau��!)1q�Gbf��n�D����ft�U����#W\���ә��=L���L��G�'UB��V�x:T�'^_���q�ӳ���[z���c�<��@�<R�\]���YS]��Ҽ�:��L���e�M�Mt9���f��qM��Fbw�^�����M��OI�J��]q�F����W=\m�b='IŬ��L�V�_��x���T��ei�'�,�m�?>��..i#F��;X��u���7�U��Et��EDtvQŋ\��y&T����Oq	��!� ���i��_�;P |�����p��	V��S~��ڨ������S
ZybĐ�i9U]�͜���mY~U�'�/�zH�|LI)t--�у��[T=�J���c�LHH)a�`�p��eb�fƚ�0���9���@��L�ۄ�|�~���f�ސ=
�'n��977��K�N�7]�
�5~�F��op�.N�W��m/ӑ�K���.����ԄT�ԙ�
��� Hd9���pi� i�f�b�­S��
�������Ĭ3VZw��������(��r�h<�G�L���͐/���8���OO��ut���c�o�;!�5�W�w��g[�@�k4�y2��⨜!V㘇��)�aL�/�M9/��M�L.�����ƌ u���i�FS���&���~ /�}�]�ٽΔ�����L����G�����?.��7��wA.� ��X����r\�]�8l�n�?����(H>���4逃J+ ��:�C�P_�3���\>3��m?E�8�b���Ҳ�~��/+���샃cV���z.�0\�4c�X˽���� �Di����΀�Yf�?4��uj�b���z7�t���MZVV��ַ��[�E�����<����1����]R��b}�G�1�ɦ�*�j�=V5>�h�/�'�gN�F�v� PT�����s}�i8y���/�\^����K蚟ZОѹ�L;�7�Xqr#sPY�)w�Nt7Kr)�Q�L�{�x�T�����P�����#��%b��E55�q�ʱ,#2�q	+7 A���X��C� ����[�����Oޯ!�����?���ݙ8������G�FC���4���G�G/'�ήhmm�%g����6)v��yI2{q~~���1&|��o��i��~:x~��%���)W�h_��>�E�g
���G>::7��S�S��+�?��1��-j�egP�z����g�w�;g׹MOϚ�ˌ���c���H}==��T1��g�i�30&n9R�=����Ӷ|�l2]�W2Sʣ��c;��դ-��.��2~P�_�E���+<��<���k�ς(��YA�jhpG�����dw{�?�lQ��&^l��e�u௠�BeZ^��e��!kuvl��sbR#o������j/�BLԇb��o�tu�W�ڼ�R�I�c������f��g��:�We06} ј�o�bzҶ�o���Fɐ=��>�QwW��wx��F�j+Ʀ��m�ϝ�~W�І���qxә*�¬����p����_xP�����RM�F�B����Q`�9���(˶���,��kh������<dt��?�̺#�����={^k�ԟ3�@R��]���&��d�w�B:�oW`�)�*'#z�ɹ�����_'k��+��j>u�Ӕ�g��7�%V�� ^p�����!�?G�.�Dl��0�X�������o0����a)�1%_S�K�-�S�ɩ5&���l8��Y�yJ���pS��p����v���"�M0ȭ��f��o� �1n
�U8&�F(����I�=o��4��諒���C+(��(�x?�Y]\h�ו"*��N�0e����C��j2J>��痣��}�O�L�K[E��-���_�}��W��3yn޾)�r�zUQ���<� >�)*��a1k��-����]sb�2�)���^_7e��v��Ot�������Vc7p�xIY~����ld�N�ͭ����է�1=������6ZC�ٟ�	 �T ���7�|�[֠"��6�ZY߽-�p��7��E�5k�6J���w�d0ǿ�ۛ��w,�r� �=��'(d�O�@���F~����]g^m%�L(�c˓�k�`ݝ���JA�n���,�6�,�D����� ]�j��K�Փ����(FQ�ޛ�;�"%���W��b�*�';Y#���=���n��G3=����'�7�6���V��cZ��h&1�+�G��>x�';�*�����NideLf(%�����5�Е>ڰ�jf���\#3n���D���͛=��Ӳ�ܪ��9=5�ΩⰘ��0�Tq�=���и�oϐ~��bE���M��@����{e�L�a�j�����@�;,�f�����ԯׯ�����?�T �
�B-�c����m���,���Y�M�d����,ѰBG|��q��%,}!�����[ki)�-�5Lz4-�]��ܼ��%/>�A��s��<	�u��<�8;*Z&�u>���6W��]�X��Z�j��u��bB���h�0!�
���?�� �6���U��C&�J�����X��!-y*���&*J��=+x�����{/�4�L(��ow@y%.�iV%Ԣ��8��D�J#�L���Gm��*��}Դu�$9�ώz.�n���]{[z\Q��G��F��5.-ed�0�9�,��-�0��k"��N|պ��s5)ļC�O���GMj�R�٘Ƴf$�%.|�Ư�����<�i��b^�\!D�:;�4n<x�d���@����_P�����1�=5PMl���U�}m4$3..'E���%'UrR��.�O�Z�MZ<���k��s�̄��w���Y�k]���5��=�yӎ�9rj���j�=�|�1�����?w�ޕ����0َ���� ��?�s�x�.j#P+��BK�0O)��\����˜�~ŀ8,�2}2�:-��S$y�ʞؗ�w�I�ͳ�:��Bi����鏺�F�L.��E���pU���j���:���v<�v�K$#&8�����cǀ��0�񝝝�úZ�Ӎ�<�R���	d����d�S;_=l5��BGUh8����I}v�#,2I慊�L�����s_̈����-�r�,��4R���Y /Uګ����������^&��@��d,1�ꋰp�Z�9PP-f���˨Y�~s�oAX3%��g�b>����K��f{�2_����j����)S��x��0!���;D ڥ�y~���>�sHO͛�&o.����ǥ�N�W��)��R��=���o͵w�Kx�,��-���<o9�o $�P������ډE�l��-��=w
�;�f��Ι2�f����'���N���->
t���ϋpi?��^���F$�e���+���r��+�?E3s:�Ap��� ���O'����� ��IG�~,����fg��`��5&4��u7�mNcJ�z�Ҕ��)qp���x���3I&3΍���},�Yw�`˛�)��?�B�ҭ�5f��Qƥ����|*��Ҹa��l�P��f�a6�f�}�+@�|?�]]-ܓ%o!ظ�p��T<�}\I��p��O��fvW���^�[�W�����DK�Lm-�k���5�̾u����3<����Ա�Ni�@C`�w�++�vY��J�䍽�r$�(��yw{�����v�`ic�T�tu��w�۔�������U%����9Bf�]k�&,%J����o6G�5�fddfe�3�5Փg6���^w=g^�ϡ�Y��k(=�ǝk�rRP���]J9����	(��p�<��E�vPW�3N�P@�ydè��W �j���ϝ1ρ- �y<0ۄ�=�R�����-I��\�����L��ƨv�����t�u�^�y�S[��M �%ffV�w%�$7�7�H7������ ��J��;��y�&-�PR2{�L:�����J[�����\h��m;?�Y1�+_���ڽ����/",,���ykܯ86�*�7@����?��y*:z;��*z�L�v���lg���5���p�y������<��@�����u��[�t�i`O��2�A��(�uW��-4��\Z���)`8֣O�����Fo��V�('���t{y�o!�/�/�(Pv�Ku�fOG9�~� �(J���w��mF62����&�>�P��ٖFFF���c��4\$oE?�g*g�O���&�ޖ��,,	;��>��PH�7N �edL��ǳG A:ޟT%���<���ln�e�mV�^�����.&��}���>��u��
/v˾[$��/X+�=���������\���ôۈ�9�ACo�W��V0Rj��=��o'y��'�|f��H�'��'�v�������ҞK+�q<�WsфxP��F�.H����E���y��{���z�����9~'����%�KN���)Ғ���h��!��,��<��,�neA�<>�c�������	ן�9NT[���#���=Q/�4Rh�����3G��kܱ������'U@����$�x#Y�U-���r�;�(�G��|�����d�5��@$�yu�o����E�~u�ct�ߧ21�&'�7����$��ݱ���F���O����/�7����n�P����|JMez�si	Ԣ���.`�Q�+#��i�Y���Oj�|����p��ۉ�dF?�y����晷��6��q6.l}���қ����؍FR�G���DR�{�A�[�&�ۦn��@�pe9ݣw H� ����=+���`�}���%��g�$~�LU�m;i�x̚���RF���qo�r���:���5r��б/��������8�Xv���f��˲xj-�7��!4v�����	M�!'�I�BM_��TY�r�R�m��7�9�7P@F���I��IA���~ϥ�ׯ�^5���T�����E����D'̓`���l��p1�Q������+7VoeS|)+{y��C2��Y���oI�I�ߤ�/��Z��^�w��@�:E����6�;=��z��1������������C�/�utt��4L;b��wGd:���A�J��I��Ԣ��f;87T���ZF�L�s�h�~ 忯t�As���4��;�ņU��\I�~���a��}*=���p_|N��5�-iö1�U<�,k?�$+��j�D�0 &�f�>�7d�1��y�( ��6`:n[&x?��w��^݊z]�6/�B�(�LB.����d(�c�Yuڨ�����!T~�r��LSu�GX�~�6����A(9��W��s�;�G��0��~���ۣ�j����(d�d��÷Ǝ���'\m�ն&�s[��/���s�Ua���ô�"����[HHP!P�߷
��?n��_R����)�g�t3�'1�������dU��z�qhO��O_�g(��(lj�1��x]DV��{��Bz��Z��{{.�E~��I	Ȟ������O�k�(s85T:�w��k<��3���J���tBp��O�@�V0��Xxb���>�I��f���v!�l��0H�Bo�&�����s/�s�K�Gg�>h�LM���J�2��T^3��F�� 0f��̘����(o��+`�_Du'h�������\B<<�ʣ�)��(g ��b�cҭ��&&'��5�˓��y ���j�VFU�����Y�F%(k_zy�x��L���G�5�1N"��%V��w*P{�T����\\�k>h�l!�_r�;�ws��<<5�]t�@Ճo�M����:=���=FGB��q�{�.�҄�G����酑�]������.��Y��w���K���!?6��~��ڨ'ZY����2�p�����3��T����~�j�+i"}w����������u�!�KLK+��L���n�4�@A#䲧��%%�=�:0G����}�G�,���yR_�S�nW$y�5O��`R[��n�h�E�c�nI'��1���f-�$Ȃpj�w��ٽ��$��ᗁy�����e�(܂ue�&�2�f�'1��)+��J��{;��Gk�w�|NO���J���.Ȋ[mN�LW�D�5+;d�{v T���@�U�,V!�I��~���H�v�/Ak������((�s�4M߰��� `����ﬁ�P�c`Yc��	�I�������w%����fdt�&9$��ш��9�1ݯ�6]��O�  5�)bvp0�SX<j����+�;��*~?��4��$��;�I�)ц�]E��u_�L�gtwf�*�n��G�I%T�U���]�n�������������R
����[[[^r�@�1<<!�oC�(לPi>f�k���δLζBmS����T��y	���_\Fկ�V��u�| �<zo�AՂ�]�Q�7ΏM�*Z�̤�j��/}�i�9�e�׼޸�%��M��M��~�<�$��ͬ�2���^�*(��¹5 ��}�Rm��%���n��c � �y_3�1�x��mn���+���[mX�q�S��$����g�"т�Na������K����:�I� �����҃(G)-�s
{��7*9��J]�2�!���Wt��c�a&P�Q��c�WMS��ݽ���C��S��9UU�Ύ��[0�,�%N�ݾZ��_U=��坑�5�+ �M�!��M���䇑�8~�df�ԗ�*裧Jc�{�5�HY\t:Z���t� :p�eႽ]�ͦrYZ&H��T��i�Gmp����_,ڰa�e�2���Nu�Q��q�J%_=��EU�\��8^�<�<�d�eH�h9 ��r�N����/��u4�hg_����^x� ,5�XV��zy���v�aC<�>9:$�6Oh����i/M�w$S%X�������?��f���f���~���x	��/'+r9G�l�T�VJʲ�7a��J%�T(\�<�}�_�ӽ���l)��Y�\l|
P��+�A�,�ְ�D	PWc�tW<��H����PGh�5A�hO^;��,��VV@�V�k��?��	�����ĥ__6���??���g���;<��
��r��6�W)����@��x��	D������M�]��_C�(���_����iy���@��6N~��yMK��`՞�5/=��I~\O[#��a0Va
���^�Y�9��uy{���a.L�o�%�~0�E���~+��gy`'��;6�i�qS�����2��D�����:�CT�$J�K��#u���K˶q�W{�][����4�aـ)?;[�ں��2@��}����띷�Դ�nc�H;1��^�L�a���ұ��w���c.K�8OC�5� �?���<o�)dh�#K�2P�f��q� u�\��ڻi����=���m��O�?:}���VW� T����w�N^��.Ϟ�k=��������	wr�'
�y��_rg���܊&#O�iW%�%���KT�a��;���qs�T��z����·Ԍǻ���	�y���I $�ҩ?�#ئzn]ů�3�����qG��v�]%�rȥ��,�[�&�������h?�����;_[�8����O��(�d�����o�-�DO2�x�ҏ*v�P��|0/#��48�@4��Vƛ�qkЋ��f���VD>m)�~L���h�E6��G�^�/?]@���ďvq$(��R?���靈���a������L�(M�����'M@�:�D���p#
Ǎl����\����'��!Q��ۇG��!x��x��K���ÇO��-�L��fJ�i�]3�"�YCf\�J`� �N��[�~I�;b��-g��t:L;�<1oh\�x*��5"g�٣�`-̗�>7���qnX��� ��gו_O�*�GgGc�����`E��
L+�>Ό!�dP|j��z��&��qj�M��A��a�9��y��rDLЬΨXD��!Pq�L������C��7��q�0`����d0�miSE�5&��p#�	�z���0u�OK�0�����z_o�i�&{�l7�N^�Y����U26W�Y�����Am������I��xkF_�ȶ_���V��5���kP.�!��|��M�س���a-"��Ի�һڭW��i��^�i�(��3eT���3-�OR�O��"X��J�c��q���U����DNN��.Z/��_5,ӧֹھ�E�xO��Yb����y��*f��.{]:;�\͂#�j�E���&qW��tz�ٱ
D�FA������.�A�ϟ�Z����UQD�����ѩ���b I��@�3��OlOw�����1�1�c���(�u{��?79q0a�fE	:0!?�������p��
���y�!�?�W�H�ߨ3Mҙ�������Q�vWn�3�Ol_I �3�-Q���v�L��T!t�#�]¸�����O�q���/�iF&-D��6�Q�9���3�@��:���>6�
Q���8/����q��!%%�~7^��<��Ng�p�Yؠ������'�1���7�i��}��B�X-�X��O�"�c�~_��?��J�!��f��Z�>	a/DM�7�(�R_�WU�R��ba�ϫfK���j�|Y�+R�!W�P���K�/hii�I�NÆ=����;�M�Ti'���-�"�	����R��3������>]r���a��厡�A��o����[��fF\�
�g3�+Pp���g�'�P�"��òg���uj�zY��L��간��vQ����Y�,Ґk#���^Ġ�� �zg9cE-�ȡ�?X�l��y~v�v�P����v"�f�����}����+��N�r~�v���,�h�Dz��(��h��odI�������u,P��U�� �{�9 ��0J�����������_�/�?��(�C����A����Ƴ�����V�ܾ-�4��?���K�L�0nxa�������(w�~�̆S�P4+��q���	#7��
_!�"V�f ު���;D��0�r��wa]1oO���&��7�����z��H~ Do�M�\������X�&�o�ܱ�D��#��\T�{��l��^����N�n�C�EIuhW�8�Т�^�@�%�>`Ȑ/�%�{��N��@�`�z�j���:��y�w'j{{;�b<rzϙi���/���F�:������z����n/�Q�<��:� �x�u�̆��F����x��[���FL��!��&����cZf �j�M˩�W�Go�-7��O�cҷ=��є�
�����?%%�%���Ǳ��5�w<VJ���H����a����m�"�NVx{u)Bl�8^�H^���p��]�r��7s�sOu	3���8t<���3��y�?�ބ� � ��h}��ޓ�Kmw���5�#aH� ���uL�+bIV$�y��$��bݑ������굯�,����_mcu��9�e�m�|��{�w[4C|!���x�����	D�'�˔d�1���Ã�$�?��չ�?�<v{42��oص�S<��з� �7��a� ����q8�����JeEE!YHj�BR�t�J3z�������.��Ѹ�̌���L?�Ϙ_A����_mf_�~�SffE^�]3����Au��)�����o�yV�>xvv���H���Z�J��:�鰎���L>�8c?�����Pt�0�[n��%$o�wֵ��k߹���?�R�;h��I��5�#��Q���9/�߯#������S���R/��Ӽ�����2ޫE��{###>�a�k��Z�eX&��o�u�t����r��Fs�t�>��ܻc�w���.�O���MIEZ �<`M7ƒ4���_���+h�:�s���_��7n�;Ӹ6����QgPZ�������w߫I��O���̖J"
]^K�Ŗ*���n|�!���;�'��9s�=8���l>.<����C�D�WF]�P6m��x�'���e�$�:��������;¥&��01B18\W�2�����?�B\i ��7�@%�v�2���ʱ-�C77����TII���qG*Gs�����_���z����펾�lJj�J�o�csQ�'�@ai��ax i����F���~��(D�{��������L�j��02`��K0�Dv�;)a+6�f?�L@}LC�A�e�uc�^�A؉��B��bG�i�l6�R'�xIdt����i�ſ��{!�rqؤJ|�9���W�H;���v��ˑ��w�/��>��\~C�T�f����<�ћ��Y�_ ���7���7n|U������4�H��}B����9��NzE�!!��x�,�84�_�
n��7�p�3o��j`�T��/�;�(|Ч�tT
��(�3U��~��GLL�1C����������;-��(Я^X��@͡�#��b/P6����֌fm��$�퍔5n�~�%~���`�>U�$j�1J�����( 6^� ؂��J�ߎ��u4R�ٗ����2?.��jwؚm�*�����Ihy,t(қ��,J�@!-�RA�K����\p�޺|ٱb>H��R���/�|�UUU�b��0�T�ommE���`���"U6���.���⛘��=�`�g������B����o��:����v�Z7lO�T��lC�q����CI���K��p�^���[��e�]?�:E�b�:n�>�Ӏ��G���B����I�=�)XnŶi	���տ~�`���=d��t�aC���|��쮽!K⸮�{�ixU%��߻g�kφ����v�j^R~�L��r��е�炇*�#3�=��aYr>��U2]�N���ݽ��W���<�n��ڮ��}��(IƯ��BϐHC��T�	�	�:�Q��y����U�[�v��v��h�4$w�����K�"�Ų�/�%q��y��j�j��������&P��s��T���{D.p�vl�� �~���.�$E����3]:)�>}V���BwJ8`��ŝ?'č�w��<����?�oI!M'G�1��NUa�`��b���]%��&�_%��<�Y��-1ih��mB����L;��C�r�~�
Q��^��_o��!�����r2�8��e�j-�~<+7 ~\{����5\�<os��F�z�c~����I���ז"����^o�(�UH��^a��[h��߹��[��Ei�}�����S�L®�֓,9(����1�XGm��fv	�`p6��El���$�t7,�k���v���d��"mhP����˧��ؾ����xD8t��w����̕1҃o[3�,Y����d!�W82=�*��o�y���#K)Jm5��3���gA sM�k!��'�U�2|�R,��������*�Sl^_�@�w3�a2�����S�Sǽ�y��f$�%��{*�����-�V�?�(=���x44��$���2,���Uvk���4���>Ӿ�f�׀��p��ثgr|̑k����BWq�7M�{u$��⑛�©�t#�3*��>�M�u�O�We�@�ܻ؈F����{�]N�&_#��S}�0��J�������gv�b�s)�5
�&jJ����S#��S	�����iP�%+�+��9�O]Fк���<z/|��<��I���glk(�=��}}^/�>?8X���6���|?��#~�4�;�Қ�� �n1�"����(����1$mz��?$���_�$�h�E`�Z����w�Kj��9���@�����_��[�2�f�)��3��öD��y��RT湹�����a�_M�Vd�8|�v�U/�����_�h��2L�i��{��h�>s���7�� Z�Pd���I�D������U��7%�:�U�� �B��=�k)�ͷc|�j������|�s#[��x�*�0�+�ya�m�BD\�~�Ӿq�$*��W�ՇҼ�?���ش���@j_sw���� ������Ώ��6ۗ	8�CJU��	�˲u�I*Ư��0jY�����F�^����<_�5�Qr�oYҲ��@$ֶ����V^I fI֨G���~_ܩ%~3'KY�0�����U_y���Jg/�k)O�Z3�� ����O/y���������x�����^���K�+}��.����zt��M��Ҙ�z;���]��C��ɭ
���޽�H�j�ڨ�T娼�e��G>�'�l��˜n`��y�@�����
u-�k���ss�E	5n��DI^�f�<���9<��T�vi
=����!�y���-
�4;�v(>im��GE�s]����4���>T�q,=H�t�4*ؙ_"/���^__�y,�����9=|�����?6o�4��]>��O�kzK�Be�U���R�$e�N�o��Xh�!�]�� �V���i��5�oT�'ݕ�g�{^����|o
$N5ݢ��.bL���>6�n��}�"��6�V�Fo�'L������H��{St�������h+WɌJ	r\mm�P
m\�F��7�2�>쭼���U�����t�aQ��~�ƥ�f	��	i�A���.	���FBI�N����;��{��k�y����̙�s�����4s,4�ӏ�1�&�mw�es�Ȕ���L�f"V;���O��\:�A�eU�����f�Ǎ����c!}��"F���)���G�t�����j>FEq�R��TuF� �/�Ê��F��F���,��c۔��Ie�$L������)���ч4�fVM������̧��Q�\c�H��ML�w���˶��*p%I���k��|��5�Y�d��}��кt4pP�Uy��|�}����z�@����k�V�zqEM���gq���3ǎ��X�lsH�[�1<̐�LN˨�c{��/�Y&i�ч�F������p����u!��s���<E�5%��� �(n�F�R����J
�t�F'=��}1������:��L�cﯻ���v�[]�E�v�d(fW�Xa^��|T9�x]�u�9TM���iH��1SkQ(X@�L�S<Xc��X��X�+R�R�����Ľ&�?#	�a�����ǻ��jȯk���7�AcҚ�:��A҉�� �Js@~N'	����B���r����Q�ˇ��� }U������-Xg����~�"t��w#��k�1��`�mN�z��Fٖ�&�.&�l��������h�����P�L���-��TLL:��B��~�F{�v��T��T�	�⒒BR<1L�u��߽{g��_Y���u���t񠗲�
�3�kI?,z�m�B8������(B���hj~�I��=$�DQ#C�y݂�|�}F��IB?�g�'�.��tt�&O<�q���x?�v�G� �l�\z�������7 q![e�Qm�"T�ׂ���>�o㫇�Z���Q��f��j�����0H��ޮwM�{jifh8�k�`)��F��;�ҟ�9ai�[q�&y�(c��Y���,h1TWw��`!�)0��(o#�h���#��>Y0�DAA��F	xH�)�5 �ӊ�,8K���@�m;��(��-���� ����C�A�陦��S<߾}[�u��_�Rz��T��:t2###���͏WKg����߳�@>�hl>�٬uR�)Z�yyVw��Rx*a%3h�4Мv��[f�l�Q�@��cck�S�/Sr$	D(!��@��44(a��_�%��� ���^�r�+��
s��\Ƃ,q�������خK�����f#����s$S���[ee\=6=���/}�U큖Y�b�K~�{O?**��М���ӗ�QM�n�b�h���!Χ���!�z5���μ�b������8�Nh�-��mЍO�T
���`��� AFV��*X��>����D�cԫ��m��y�6��.0��a�|�����v�
^������pP߆��&���a���u����l�q�{��J�@��\q[������[rr㝻�k� ��'��:JTD琱)5�yf�Ost�t�C쌟�E!�jk��~;.���|��eљ}�rr�:D�?���t�����:\�����ǅ5~��ˣe1h��+vȮ��x�eז��oR�ˎ�p��Aڂ�IXj��.Ϛ�TRa/@q�"����0� �ۢ��xM->VZ�ZQ��o���X
�+E�?�2������V��}&���G�9�{����fn�����3� ��Q��t
!ˉD��#o1P��*� $��$Z�/��LHL�f���2���b��4�/m��gT�&�/�=t'鐲��Y0�3��iw���Vi
zϐ��7G~��;�x��=�=���n�-�#���Q#�0�VY���`��B�������"�x9AUt���d����#��F)-�2���<G�W�n/?U��5.�X�����Y3�^B0��s�8>�iF�=āo��{E��1���*���"k�)?Y�`������n�1qiā����	��֭��U��Z������~�Ȉb��Ղ��˖�I�F3�b���HEʙJ�|����������1Tx@������ Q�!"c)���2�Ȍ�P&iK�C8Ù����P[�W��C�橪�ZXٲC��%t�KT�Zԓ��,���t���������YCKk�l� ��9�1��tΉʱB���}�U�L0���=��j lf���I�	�ӡ_�$�mmG�'����ń�1Q�����st�X�Q0��u7�X���#](�� �w\�sqq���=�^/;��s�T�7mX��,��/ݗ.K��=yi���`~$,%�IYI�����H?��0&&�Ii��n�j�2��[ۦ��u�I���Lي6F����Ҙ���N:#{E���:��*�+J��Y�y���{�t��`���l�	'��X�e}o�Q�BE��3�R���fada	΃�F��M���8TY�	"�o�6����U�d�,;�C�\;�5K���b/?�עnc��.�m/�s�������/��?G=�~��E�bugPSm5��H;��e{��9��c1
�*�5�̜ET\<�T?�J��p�E]�wG�V`08A�6�:����v`��^i��dʈ#�b?�Q^��^����u��������՟��.����7X�X��� '�z�T�f`vMZ!�=*-Ny�k�_�i�]�/r�pG���z�!�˘N`����)2Z�Nٓe Տ��||��^�ai�����0��>�����;v-ޥ�H!��A���vq����#L2{�b �2<\i#��zt-���̉��*K��A���n-F�i�1Pn�:���>����8�+j�ciσLz�fdn����+���59��Zϖ�b��c��C#���J�1�L�Iv}B��Y>�7��y� }�Q��L���v�N�������n��I����ޚ'�S�-�4 �h��
��:�4v���$��d�7�{���9����U���]͡O(��?B��g`��a�ڄj�k}w(R)���@�$k[@e-/�ioM�b�` #�P��\=��v)���O��T��5A8�=�K����>,�{M�{��ὴхMnfu��������.J�$}�v~�!��!�ąt����U?��@����������;��w�X��W[�����~��rty�����o
q_������������P�����(zh����u�Ģ�2��>_s����i�@b��}��sbc-�8�0�xuw9�˃���<3��4ނ����+��}��-��t�w�X���._�x��X:�<	Й����Xj���
x�3R�?��u��#%�e?f����oĠ�� �h����o���gP�i ��늚�JK����ߦKY�c��:O�_DEس��ɬ�_����מ�'��ѡoRn�E�F���ȴY�-V�t_ȡCW`�_�~���<^�b�c�0��1Ul���$��''<��£5�)\�ƿ�eZ�J�2���ōj=^j�����E���'���W)9���w=�PJfL �M^���m����'3]�Ű�������Ix�l��]��q��Lx�u�3ж�r���}"H��зn�|��H��SG>\i�c�߹��r�nں���s}th&�!X�Ppj�lЊ8s�[Naؙ�,pB}MnV��hYo���S�~T�n�:��G�e�g��,��2Z��~鱤\fr�!A�T"_�Ү��}��m38?Ә-|[���7/KI� H�G9ߩ��/$�r�8$���1M��W�0�� �C�M��$8.;������$QwM�l�XAY)� �R�!عm�k9hJǟ1�V\� ���,K��v��������w
$�@��P����O��j��jfk=����oE���Q��Q}�t`�*�����kf�+�v��U���%j����� �nk]���>3���G7;�a��������#�É1b:J����X����V ZZ*����C��;I;�(�rm:�輟�ip�'u���lٟ�rh�=�o��ί��f籌b�_������̻���s�Ǝ��p��� �4�ȑ�n��O����/���읯1~Ƞ�n%(�>B*�[�������&��n�ۍ!���x�O�e��L�G3b�1K�J�n� Ω�����(����Э��<�R`#���<F��������i~tp��~�\_�E�Z.��+��܇��:9�����d[&��Y�����l��&D'1��4���0x������n�9������W�񯜢U���R2�}7�m�{9��[�qU��h��րˍ ��Ͼ~̾b_ê`Y��m�mN��	���u/��w����&zN �0�+��IAr����ƾ�Ц���ȷ�uM�J�e�����
��Zܵ�I�E�T��w�Ji�Qq���d.�;��*�1Ȕ�Q��0Hm���㔱�M�pk�DR^�/�%@9t�c�.�4�瑭��jh�zkR�]��׷�dnv�d�H	.�Vݷp�����7v0h����������/O��۰~5�q��f�85D^�/��D!�/͘b%���l�;��T�D
�i��	�������qCZZ���m��_�2�� ��g���9u"�-�ɶe���x��qTs��騋�Pa����ʕ��m0.P�HC�������D�=�Ô��]׉3%��n����nDTTTQ���l^c#�r1�������O=,�f���y�Ae���廟��� Qqqj4\
g�V���23W6@� ��4\��,�>���w����0�'䠞��K@<��4"�E�e�
�%7ACt�C~�3 �աs��ds���e�����f��������՚�����}���>+qP�S��K&�� z��v;���_���!��8�(�����C�_�nj���y��l�<t��ɤi)Ѧ�v���r� k3���J�L���3�f���Z�$���$ɿ<�� I�@�c���J�4`��(t(l�ȃH���2��O�o�ҳ'�%���g��<���������5>�]���!<��Z@F�w~f�hZq%�^2�N`�tYZ�1H_S�����٬�mMw˭�Y�!R���-�ۖleѡj����(233p�������%OJ���̉��P<y������_�Ua�r�L��V�y�~o\�����"�c�ҳ__(N��=�d�V����^�1���e`,`w{�7�p0e�/,�*c�Zik�t���]nm<,u��ǩ)G$����W��N��`�Wc��]w(1e
�����^����>��'KM��Z̫�&�vۛ��YX�20ì���6�#9��T�Dt�ΑP/*>6�57C `�|�k:%����K�YO��i�ܽ�a6O�֥[gOLm_x&�.���rx�W@�`�a�L�8���������+LT͇���������RSO�w�,s]��"����x�q�V��/��6oζ��[��%���~1d�@�͛��s$DD�#��7��8~���U���?|Ҧtj��}�O��|XA�Ԉ�Sm�$��2}gKA�x�τ�禵$|5�n�g�w��'XJ[��U�NM5�c���y����Zzzؠ�ϵ����4���R��������۾��A�?�dM�x�d�2�S�*��3u�Uߓ�o��;�a���]s߼'Xl27ZZZ����z"����}��&"-hӜs��ꏵ�h�A\���q	��>SJ{���K*�]��/��N��uGY���T�7�s�G�Q����Sm]�P��ךv�����X[��~���Y<1Bbx�y ��H�2�:fz����+������8��r��>Ys+)�k�V�ja��Y��� ������$���{�*��$�>������55m��(�Lo��ώ�fc�m���Rc������AZб��t���'�1��?=���81�}Dq�wN/H�fB#fU�ޯ�gڮx�xqL���GQ�ⱀQã/j�Ա4<���EV�'�,/�������KBL��!�4���#g>1?�x�������!��J֩����Qa�͐U�������]�gA��C�o))/���-�<���� �Ib�����E�&��hW.(�)&!�\�1�^��T�������B�{r�����T�����5~�9!U,1K�qg�t�X�9����՟�KIl�ͽl�?�A%��l���㤦)���&����BG\�H��Q�9��S"��1G�<�a@W�N�x���5(~��"�	���]�3Q��t�R����&|s4˴6꧔���3���������jPU���e���|��5k�j �*�:����5�R'k��#�.π��)�B4X�͕�g��׻���H0�i�*B��*���ilPmշe>�I����3Ass�A�x�`�@��}��d��IT��`��Ѹ���׆G����G�牉p�ˮ�2��������d�G*�9&�r�W��\@�=�.<D�֣
��-8h{}a�S�ţ��' q9�	��حu���nI�����g�Yn�[j���b�}�9��+�rV��wo�N:���b� g3���d*Y���	J�y�)Lcq$�7�[0jZڸ���#O~f�}#�����1�trA���o)i�MM3�ڧ�`��oefOJS�]�Gs�����sd�W��d���w�8y�E�n��]�{4���"�R�p�⇽��O����zS@
��	j\�������;8QV��%���K6>�F�TJ�}�ev�[K��T"`��*��.��;����z��+�����ׂ�E�`�&�~�q���K'�%(�-�t-`k��C$�?��>l���t��N���T�)6 ����9w��(L�;���ݣ�¬��}�D
�k)����#2�^l�}7Y0]i4�b�d��u�p������K�;�e�r��DiS
��3�#֑�)�=yAK���z$k�@��dKQ帥m�����}Z�xkAO��#�2!�8���?�;ׁY:�Nԩ2�<t��_l.�����[�b�Y ��>�K�ᗔ]o$*����Id���@�z1,�%&��m�K֊lp#�A)=�7����m�����`���K-�g/Vj�ط����DUӼ�G��x��Z+����U�rW�G�\ML�\ە樼$+l%�J��/�]Oly���|\⑄A�rq$v�L(z/r�����NPi�hIy��f4C�?w��j� ^Q���8�imyO��]N���m�*RS�NÀ����5��Ǵ���j�)������_9u�7��y�)9����#�tٯ�'=U��ѡ��JK9�Pꓒƕ�K������;�Mu[�� Ipڢ��ju�ih��O�C��޾U/�2�)�Qn��g?�jY�?{�% �$�;��	�N���F��K#l�.�k�����J���?�'���iݏ���Q����!�.ꟸ��`Ć�w
�P&X�3�f��0������@�F!�7�����}��ĉ�9��Ըa�]d�]�4�8�mw�4�&5���2p���:'��][�1����_~�� N�I忰(JC�	�`�e+�����F�,��٩ؗ=�r�xZ}�=N�֞�� �� ���y�gr�j�@PY?"𣩉���q@(1bY��n/��چ���Kr�Bt�8��U�,I,�GJJ���4>�^���U����,'�A���L��ZB����a��ųO<�;��Jؓ���\`N���魷R�P����y�|И~����i������������~Is�aʰZ.�g��Y�ǂ�_��p7!���gnf��c
������$�o��U��6�_c	��\�1`keTi�k��8�+p"	 ���K�����rZ9#	��W�~E;��yb�����NN�~�{�Yru>�n_�7�X����<C���u^�(�TyG><��3�X�1]�-��9��s�kM�p��l������JU���ތ�1��%h�A�Qc��O�U���l�nY�GW��Fٓ�=���I��ő���q�_.T*We�X�U���3���[����݅��[��n��U�1��� $HƊ1��m/�U���[0�Ę!%Fz����'m�{vQqY��֧쥍�0a� �}�H���E#*t�I�B���͎S����y��|�����@��m�?!���飨��h %��z�����Q)9������{ ����D�#������K3��m��[�yP�*�RP�*רn)G�н��~�k��w���G���iWV�?�@�q�8����7+N�S,9t�}�����KR̐uW���;F��"�SO���2YF�	e������Z���I�È)�XٰOU˘�xT������Z��M��S���}��F	ӂq�6�C��[�5#�(n,��U��DR��d8�
�����	�E��
�Ķf��H�q�j]V���'խ���\hRRSszf�o�z�[�ܜ��]1�<�r���Ns����Ў���P�(�`
�'��YZ�WYI�$A#�} ��$I�U��fy.�7�	T$�����:?9��*�F�wIt|(�FM'a�Q0�2�����<��o�(V�N�
~��\t�q�	b~�{�3���0_XP
]^���y��� q
n�K45,�*��m;��`��UJ���7�Hh�,�z��Gy@E���	���(�q�~ۦ�I �T>��Yo(�e�y��I��~�#M�3>2Be�kZ�j+7�Ɍ��/��	)%� 0�H��M��¦F��B�w��M�Ne72g&c[�Mm��+���i��8d�c严o#G�(Yҟ�����ʾMU���|���O���k8-�pG��885D�t��p�Kt(]��5w����|�N{l�e�O	���gUF*YI�A��T}gO�b�8h�e�{ v��W�ң_��3F��*�I冾>rVO��V�"��W������U>�De�`�*8�҅�\��|%�j��F��bGa����4d�q�,�\"Yqd}�����]b��^"Ԯ�b����A4�ި5R��Ku0�4�9��*ڤ͢�2�Pʊ��xT��A�^5�ҭs�w����s�<����.ʩӌȓP�V�c/��EN�b�@�K��}��8ʌn�` TR��7��
@��.F�[�~���>���J�U��*'--
:Qe��P���PI+�J�n/@�#K�(g��{S]��~�#4����a���a/T^�k��,�I���^��񍷤ƌ���N���������[�H(-w���)���H��ѳw97zڀ�_m�ƣ��Kê����6iթW�iq�G��Rc�2	��˦6�Nht�/GoZ��%�5nZRU�_�8�Cۤf-9��=�.\��)[ߓ�c�j|�.XE�y^w���RRX���ǜ ��-�뇈��s��dAǖ	�a|=�[Pf�����vT�QX�/,-�ˉ��=n�(EG��<WA7`��u�*�e%	��ꖕ���,�8��4����UnthQ��96�$9 �#7�C��0��wM���/m6R���R;�|��8SW�E�������?H�v.+,Q��{)a����k��m^���U}G��r��(j�9j�ÆZM�]ty�kj��y'�N2�K�җ��Ḭ��$��3q&��o%� � �8l�[�*Q.�@ip�)jn{���a�l��E�{�,��]�FQ�k�>*��� �D���e����w�h�[l���>ۓ���W-lz|.<��QMO')X�������y-���cY�k�˧�������wp�K:㨤J�g����Z�,���L����s!�j�M��L��Rb��l]ޜNQ�w��}���F�K��>�Eʽncs���7뛰�옖\��[��1��6E�g�I�����(�̐�F��]kk��ٶ��УH���9��Y�0K�&tM�؄L���ATMhc%YWZeD��8\��6�yP�Ҋ����E!���f:?o��{u��C�cd$��>�y���A�H��j�E��a͠�AES/��+�V�g� c�b��cXF�O��b����L�d�n�bB���]��t�/�N��Q�u���	�c�@'��w��<cgY{�㐠>�b�O����������ei�{;q�9�T;��t=�O�ͷ�NƇ�Tm���Ţ��z���%%%�@49��T����Ջ{��9=/>��lF���~.�(T+�x��:qP��a�� o$ё��i�e[Iz�l��2B`=���h� `Q����V��L�Ԍ%~l�)��������4�4�l����z���!$��a�p��՟)���v�����m[}/�mZ�;}�m����gL BΌ���K�m�ZeQ־�T@�-m��K~rw����غA\�Չ*1�K>M)�����ش�W�o���$��ǲ"��
wWJH�|^�=�f�u��(����"0R����X-��Uy~ �;x�U�5�����ׯO��O�n��SLa�������J�����K�e�*�T�bf}���������آ���>�s�����~/��'��4�[0�U(�����Wn�-xI��Uy?�2���GF�l�//B���K�����C�Õ��Q��Aj?���+2� �e��٥J���O�x�\�(K+��I����_�wL��J喯j{���KaP���K>�/�1`䤒,�C��@�b-�8��K�;��1y�Z��T��Ƒq�gU3���~l�I�?�!Ǡ���6�1�A}����[T����{�a����-&"�u^oe�z�0`2�{�`��73���>Tß~.��="��V���w�#i���%�_�ܘrX�PT��":O�)��vQ��Lw�Qĳ�PpX�%aOQ椤����Hl���t,CP�y��H������|0�#���R"e��*g����3EL�W�w֟5���)[MV��ߊ�>��팫~��4�����B���ִ陂]�j�4z�H���ycE��v���X�����ʂ�+�T���szN81��^'$��n�P�!9�?@�	��tB�H�8��g�B�z��f�-��4��G��X&dy;4�ٸ�΁{ A�>KF�NxQ�]ڨaN�+@Lo�����G�u���M7�Mb^P�
K�m'} �4��������c��~���V(�zѺ���"��y- ����6���v�DKiE�����q'X�V�h��M�k��fg�VOEx"�!L����Fcly󡹸+%kp�s1Aasb�"�K-V�.|�r��$;�V�����>��/1�y/���jcR����|XE_�������+��H8��>���A3LD��9ϧ���®-I��+:[��Ʂ��Ɩ��6�����6���^�T6;�1I0�^���te�U���q�8��g���ݿ�Z�~~����]�NyŲ_D�� K��4A�1�cW��0W%Η@�K�t�8���n5����C��娀�Ap<؞M�i��؛2���������,u����~��d��<喳E#'�x��˚�'Et�2ʀ���0����z�
[�Y*P���қ�y�
l3�mþ�6�ݸ�Z���r4.�i(�7`�2�;���~�:K?X�#�ĳU�F&(���w�/+}�z����:������SkV�Ⱥ�?ɉ����A@$1��7ާ��a��y��N�zC�f������"(mWk�\N�Rr	�GG�m��*
zm��o���	�Ԡ�p��#%h$�ȸ�m��C�!�7���A�B�� �T�`�awG*�u�\[�/W7FϨh���MǬ&���BG�>����X���`�qI��K������X��'Af'[����l���iW��]i���-����ɐ�G�����bK�9��y�]��q��m����W`dV�Z�Ray7���[�C���W\�Q�083&�6X<-���c�<J
�i��˾0ud��]�U�3w��M��;�־[�W_4 ���:E����@���"IlZ��؟���o{��]*T��`?N��Q(�l{Ja^���H�������-7�uIP�F���_��]�����C&8���hFȋ��Z4��)ȄN��D1Nk�)�0�#YR����s�փ�tPD� 9��� __���E'��4B{"4:�O�&
��Y{("�4�u$��3��۬̎���j�&���:1�%[\�H-�;|v��S�챗Ĭ��:�w_noA�G �tQ�_DF�	dyA�2�%CD �eZ	��/O%�X�us*B&Q�1�6��XĢ2Yg��B��df��*�-�X��CA,�gm5�X�����"��U���áS�Lǧ[ҹ`����'ɐ������(q�a���Y�`���q����׍�hS�`;�G�HPۜ�A�d��hr�R�nA<=� �"��$N�zxH��K|�o��,)�=Qik�MТ$C�0$�CV�s�Х��]�u�'�sw*�����2���&��W ��8-Fs~1w�uc��2�w�Q��������!�)I������9�%ƜH7�C.� ���{���y��o���e�-.Js�!���)�4� ޒ����*�V�;i�������g�~�(�z5�mZr� d�]���A��;3�^��d��I��&��4S�<��,���0ʕ)nW�K����GKYҐ����w���h�Ŵ��^��8�2V�I��R������Z!��hI�j?Āϴ�/��[�1|boa�74���t0F&[lg�Rސ�����L �	b���$�@��c�"����t2a�tP�� �H5X�L�u֓7��J��w��J�aǑ�n��I� ���i4�qfLK��y����ŏ����_�D�~d�M���zUr��4Ʀrj:���z9��S�t���I�p̷����/���X��f�|��˱���g�u�bM�"@��{�#݇u8�ƳD�7B�u�r�nC�����5o�G!rM��h�.��w�fp�C�|�j�?�
H�a~����'��LX�i�����&;n1�����pU�2��0G�r��$�A3���P��߷ȹ�����0;�S�r>�XŦ/@�a�|�BO��Flt#M����|�y����� ���n���,-�6�����[1�>w�ws]��>n8��^�s2]�ek^_�Ǐmzub��u�s��l�j,t�Ўy���7E0'0`=%�Rz�0M[!i�<҅��[!���<�Ὸ���B�M��9�9�dl$\�WG/��S^����^q虚e �{PbNȨ�$x/���ް����t��T{�[�<2�of8��cp�t���bC������+N�9H�.��P��r��jg���6��^�vT,�n�ɫLom�}��}P�߂��r��g<"<��7#@�7݄򂦜	�$�������Q�u�{_���w
J��Vr�,g���nj�����_^}}	�ș^q Oo���M4��H-HP ��Q��<�ߎ
�B��N�c�Mk�K�[p����x��qfmZ����A��T�Fw R�ΧO�۹aT��p����bCCC�Ӯk�S�ب�-Zw���ߡ��N�ꃤ}eo�F]��x�<K�(;n|�ar��ˡh��w3t�cx�Y%ky�kZ�~~B�Ba}�71Q ����N�������=�"Z��>UX��(��$]��`a�����$����
:���$r�7���m�Y���.�G�3�h���XJ�b +
{&o�pv��7�T��q�Ó���ȡ�#�e.�Rj�A�ߩ�|��p��H(��|����i-654��b ��~"BX}�>׼]�ĥXd-rX��7X�bglx��_s�<�@����O{�O��ۈ�}�Hٚ�/N������44�CH��Sc���1�<�F�(�g6�8W�:q*HL�!r�kd��zo \�m2�]|�k�� ����n�G�|�η\��e5��_��U�L���̟Ӕp#��8.6Ǭ2D<� �Wm܇��%����J�.L-��b�,f:�VS#�Jy�Еut�:&�?����|\�g�XP��B�Ӝ!������c��L�w�Q����jsZ�;�K�qv���@�3�K�i����$��hj��>�dHN��*��K�pT:��c�e*�%`H�,3B+�0&�O�b��^�u=6����hG��p�R�+�kPx�����\� O�˜�;���#"��L|;�I�[r�9���3��sR=qx��aA؊=ji����퀞b���[67���A���`-�"/�5�d������e��'���:Ҽ�f��}�jW/M�(C�%#C��<�nh�����j	�H��Mn�e���p%���Bg]'x��eH�o�Vٸw��P�I���:�C9�.%UUs�b���Yڗ/����q��"#^�SJ(@�3���^A���ș�uI�#V�ʌ[�md"��"%ao��튻ꦧu�E�1t�(4wF~��h��tV@���@��@��fff{������l�{�r_8��I��b�{T�;���Q�J�wqe�
����%���~�{&RC�<� QB,��AU�U`s)�Y�.r¤{�p-X.��Gk�= Ơ8���!����&�_Xމ/�嫭��F�2W#������7("J��q����芧&JPq8|�ؕB��d��t��#�KM�:����e��>���@�����:N<�^n#�/�M��3T��D�k�閑��9a�&z9T���tސG�
�{ٙ����-1qe��[�UR¹:^�'`�,:�8��z�b;����y�JAm�9���ɗ5����`w��k��O�l��h��ս�p�r��և�>+2�Y10V��0u��Jz�w v���*
��8P��y�z0I�,c���@�sߊ%���_��CO3�2ʒ���ct,���d�;@����%Z�z��}r��o�X�@'w��)�������������\Yq�������_W�l���qٔė=����+(�T����u��_�:�/B���sҘZ�N���zu	\N5K6짤R��妄8#`Mɥ��0w0��*�1��<��щ�ť����Ї���N1�/-�������`�t���+�CyG�6Hޯ��Ӝ���E�˻�g�Fݠe�aV����4-�Eu�#N>�P������O�_=���(U��o'�Pԟ���lP6'�?~Չ�!�[~%�:����Ԅ#��]T�9��m���B�4����ΓT��F�_��w6�P�g�f������� ��]� l���(����­?��2����/D�|Cœ|�겍gJ5�l���,�c�����/~� ��7��Pz�T�v����A�㸛�&,��%�5�e�hy:3a�c�Ӗ?#y�!oKxZ�%���V%��9|��l���_u@�!�Z��?�M|�YYqO,�/�Kf�w�Ng�Q{u�̦���.3M�w2�vR���ɇ׽=>@�DpA(�o6�8��e������֍�����w_q��F����ys�+�!�	w\ج�j^?`�����j���AT^�5L��&
å콻<�?ڙ��t�~X3�<E������t)ע2M���	s��`���d4�J�ޯտ��̻��ܣ���!N]��)^�)2"A�ˏ=��%��^����Qu��V�lN^vb��͘�B M{=��j�����A����Zp�YXҀ�]����������*�V#>�u%%%�����RK�8"2Ҹ�wz�ܳ�y7����qx�"��y�m�g���^ c#��lC)t����|��}��n���ښ�u)Y�Ӟ�͝S�S���������8�r�x����B/P�P��y�$-����ǖ!���
���v&�h�EA�SG�1���5�qZџ�H����V�/|��M�N�;�[o�f��WJ�R���')��|=M�h�E]nc#���!��?��A#��\��N�,��jT���œ�g�X�+��z>�3��5#c�xb�ĵL���b��i��v��i,6�I�6�#
�/��f+�I�I�ɕ�~���~"�i,���&C�T�X)h���q��@��M�e�۪r%K��jn����fB7��E����.N ���YԾ�]q]��߳�� ������U<�����f+>���6��`߃B"A(ﭴ�d�=yLOO��b-�%t����_��E�Z�M�lA��.�UOF��+���b4e�2�?�!������BC_�Rn��v3K�]#�m+[D�Z�R��kӨ��Me�]iڽ�L*c���Eέ�ȳ-~���>px���q#@���fW2$�z�q=Ծy��~8l�����ˏ� jO�����D��-⏣Ʃ,`�b-�Z��:t����<B�Q��YiǙ���F���ѱF�r|/D����ї��DS�d��Tؒr��
��kY�e��ᾩ�O�p?��"��&=�c=��5`JSw"�������pē��}�v�H6����٢�s����|��˲�Tc�1����9���J|(�>�.9�y��,=�9�C866����nd�ja��!�{�1�S@������Y�����q�����EihO޺�֏F�2����3Y
�W����NVn��1�ҽ,��:�c�*F,�t��γ��ϟ谡��A��Q�5YR�82wH�o�(��<|(�s�Q�v_tiW�L]Y|&"f����@�a���~-୑��N���А�LH#��m�8�l�A9��ٽ�p@;UڬrF��H��j�1۽ZXϢ����uІ���bK�F�1:�!��>|WW�N����K�%�������QQ~��C��Р(��R�t#��C������ ��� �]Cw��<����k�k����ܳ�����pX�Պ_���d9�yu�J �bo�5"��Ṽ�c~��N����*!��ݴ(m�ɐ���`�������y���c~��)[��̳����~����㳇��w�
&�++yRT��O������@u���ט��7�Egg����Ix��/��Zy_�b��� �M!����PPֲ5U!+3�B�V�?�E3'�1%�	\���ƅ�18;hJ�;���3!!�	�fq��%�F}{k�7�p��-R�hT�4]=EFH݇ܯ'Sc��D����W]�v%��{⇆Gk��>�s����1$��aA@��9L��\�F1�	��v��'�567�ͣ`��c^y9�s�H���s�i�&x���&�����}�z�����S��[��|�O�ۜ��8<��i��-�l�}�/UQ�R���0/�%�EEy�xW��m����B4*7�pLa�iDZ��4+��1�a��F�����w~d�x��?��τ�4�[j̻D��Sn}(�>3%�@#E�zt�rH_�����5�0��4�:@����uo����=��QPS���~����<���d�Y���Y��%SRR�|��lу�:U��4��jE9w���v8	���Tf��F��Lqbô�X�g���Z��&k�]���ر��M5��+���De��פ�����R����[q�Z�g��^W(��|4*�!z���Lk�:�㤪b���Έ�+��|��D&�r0�<R�Em&�%��w��7O�"RL��E�q�v�z"�����ҧ.;�:x�� ��x�˩a�s��є�c��&7����Rh�2s4���}{?�%� $UT�GW�(��l:qq���7<|����@�Ԟ���	�&Oi����Ү
����\¦
v�\�O�D�ى�ִ����1��w��.��p/�"pS�F�Z1��46�F����w��p�;QTǜ/�I/h^���#���m��4х?�&��/9�Z�w�sxt	1�[#��"��W��c�W2`����ō��x������>o15]���N C�3�����	�����{|���<��U��Ff�,��5�4߾�x|�Ā���"MX����������њ�uׯ:��7" ~é�A�Ղ)���S�ք�c��T{��J�ة�>?\���џ�XV�C�c��ڗ4����}ߚČ��� ������Ƹ)d�-��v�h�O��DZI#�Vz<��&���8���|���u�ω� %����e~���˕>ƴ�ݒ�荁�ͷ�*Is" U��<9==`| �}�����-�'����M��*%�>ԗ�>�|0M>\Gfޔ�j�q*O�9��EA��֊����猸~S���n���0�"]����%G&��r����z1�he��]徝�t��3�����4����QXiwX��U�L�=�!��r� �ƊI1��G*��������_|�����b��=ô�ӜN���(��)g�3��S�,�]қ�n�oGt����a��<�؁���\pd(�2�t��ư����'
�F��E���ru-�p�"��V�b�I�"��jL���%����E��r��z�ׯ���J]���|n阠y��DR#I7��`������	udW|[�����E-dE�viO��g�_�/�l��~r5Т&��J�
�}��l��ŹJ���$��c���b�|4m����p��a@�$����W�ƒ����#�������,~6~�)r����E���T�����N�"^DWPc��Hm��!PZ����cr:�֓�Mh>t,֨J�'���ye���?킓�He�t9�|o��O��T��&f�c�sk�0N��jKQZP4�C"K+���TLE�o�������{��аط��*������/�r��o/A�V
?���l"��U��������n���;=�jQ�5P߯���5�[��?󢣕`�����;;aE.�����������R	�ϔ�gq���'6?/��ʾ�a��	���rAޑ7){����'��y?���?v���s�#��@@:�����[c��"@yu�[�iэc�_E%�dͳ6������X��xqu���{q�#|�Hl������x4S�߿�ۮ����5�=�7M���imݎ��'�a;|�E�I�<����t�>��?cʻ��X�&����d���wI��2���uH���p�;oM�9���i�,b��K�����@����âV�ur@ʢ/��O3d��S��+'-��'�4�L����6�,h��s���zh�/K�j�i���ݭݩ
�T:��4:��Q���H	i�N�z[�we1PU�*��J��m� �
gCw����Af�K���K��\�?MA�Aoi�ۆ��"���r8s3�|��T���� � ��O�/�f��==`|o/~��RDН�h`�i�g�y$ ���}�il�w��ҟn��yͮbu�d+�[^���/g����v6Q[�l�`w�dUXC]���پJ�Φ�=��?f���Z�䒷��]���e05�K	F�5W��)�嵭
��I�*�)�.+�U�Υ2��.�K1_!?�س�9ۆ	8Ѣ��7����÷_��<��|>�L���,A��wHw�s3�(�Ė���c��v(��d�Fo�Ћ�v����Ϭ%�Q��Hl��\�!-=oN���J˸�zB0U��B��-��7$ ��L�8����zn-'qކ+p3:�8��_&��m��p:.��{�ne-���Ԭc$G�F�H�OVV۪S�CM&�^��ۣ�����_��M`��ϣ�$9ٍK��/�|^"n��?bM��"=�3C1�<�Nj�",Ou=9����?,��T1�Py�&�'���ݸ�i��H���)*��ܧ1��P����oy���l�ao�*e���^�礏��_�Z��$�H���A����{V�T�Y(�b��w�޹E�+&�����#�߳梩�φ��Jd�}+����
�Nbm:�w�7O���PWK�|���i������N#Do:�]�ԁ���+�]6�b����Y���i�?R^�}�o-j�}}��Q-��8?st���5(���x��d*)���.~�v�2P�PV]�k�.��E����c�G�"�"��-��r �����nBr�I+K����獠n���sE {�.�!'�I��(H+E�Y�;����^"�
o�s��]<�֒(�7&a�厅9�����K�����.��Ǡ��`�]j�|�#��;��ϩ�!�&ާQ�8)s�@�0�AO��MQm}u)KI=�v�j���/E�ԁ�O-tD�s�XW-c��q:���w��N��I"&z��&Z}9#����l���4G�0.��,!�.����>��w7t޾� _c�ƪrv.����)�X���s�'�W~�*�X=��aΥ�x�k�|p�f�g�b�?��uF��
���"���ѬEq�>�k2Jȧ���Ң���T��xc��F���qC���^��H��ɺc��R3�[�y��j! $ՖŢ�o���9E��x ��;wЙx��t�+�q��ky�*��S������P�J�	��\�hb�\.�}�9v(SU����9e��T_H�0h+���8�� )p�'�N���<XgA�<�G���f�y�G�+�����L��Ѐ�U��|��B�K�������ǚ�+Ea��;/�Q��7��]9���Td�,�κ�;NL+�J�� �n��n>���V�!7%� ��c��@&w��8�o��/7��^���A�t��T���c�!"n�0�yzuDuV|h���?2��i�������)��Lbo��27`<�ld�0 t��� �!Ԥ����i�/�8)�h�ڤ��Lsr�a~p�XfĘ՛S
"����U����I?3���O�8�o���Z<�O�5B��^<����9G�ܳ��*jےD-h� �4�'����!�^��,�A���r�'ܜ�S?�e����Z2J���z����ғ�a����qُK���΅�D�����?�VK�߰G(�����~�F��g�/��z���������rI$�a@���j%��BQWO1Է�2�羼j �����R�q��#��z�%d|��Ds�V�$��a�_�8T��s����	LZ����^��6�B����n(��iI\��*�� ^�t3��.�j��}z����/�o)ymV�������˔��:�T�M��ct2�Y.LI��BD�:���Q��Ϣ	����}#�����{E�u��3]�!ο~^�
�@E����J�rG$��P;Ɯ�C�?݉A��P�&v�A�����# ��`�S�b6`a����\�wY989:!C<�\0TO� 6��٩�>���w~��*��ý�L�!��P)>���f�qP��(�zz2�Db�n�F�D/�MH�%ΣX*�ͥh�&?G������G,;��������^s�K
��{e�K���'�D��v��y�Sc���/ys����>Z��B��1�6��M:o���ӗ^W_\��e�Ŋ[C�~
�ϟ0�I����OO*�o]��vB��;5TN��A�����5��ܜC��TJ����iu��Α�]�F�T�1�y�Ez~��H�b$�*EA�z��Z�~ԟ7�RZ�T��O{I�iJ�`R'��Lb��S��*�v�CF%����Uo�R�N�޸򑵶K]�:\�}{�H����(�Y�>��k��DKݟ���Hδg��I^�_-���Mc%n�������ܿ��؍���F��g��k��5U�&�|JI>����T�����(Z�ً�@���%�$�=-	J�[Ny(|t}Ap(����y�9�P�D�/�M���_��{Ѻ�����!�K� ���9g�FRq�h�F`�,*��Y��f�9�T��eߪ��~[|N��t�9�&@�
X*���*ʺ���	�
�.��!� ��^<v�łn�/G��(�e��%�3D����3Yq�nU���T�3����X?jPV�ap��ǿ�]�Y�)ԁ,�O
T�v~aI`xi�W��tR��]kS��K�[M�ɅmxFH�^6����+j�l��@p��Rڐs������c=�lD�dS��-��9��ĉ 8���R��&�|�_���<�oJ.���jr�]GI�;�Ⱥ	�0Ʉ����:�R6����<ƅ�7a�]���B�����<�&��z�V8�xY����l�2O���u�_��F��[]CZ��/c�LY�8��	�D�3���{;����`�� ^=�{��Zgp��uoӈ4�`�3=��&t���x<��F��6ә��<&Λ�Zԉ7��&��B��B���M�G��b�ݿ4����Ua�m�$��J�yw����53F�CC`fdAR��1�\߂+ITG�39��|�R��S���� E���M�Y[<���_�	PAs�9�B�8��%���[\~$����n)	8D�_��2��	�*ʷΥ
>�܈*A������e�[IC����,�B�����&�������i>M�Jv?m�!��<�$(GO�e���E��-����{���}��8��8DE���D]���1m��S$�è�A��r��
H!��dt�{��5*��T��+�AQ9�G刿��o!��q��������k�H���w^¤�E��p���������Qݰ�ϝ��Ga��s��c\_+�
���(��Tl��=$LX�r|���p�|�!>Hd%�c�ns��2�I����h�%t;
�6N�My��Q8*fC��6P%|G���0_�͟eq�,�T?
�~V�dECJԟǅ0I`��(!晱�N�cS,��u��+�	��q� �v������Y���I��Ѕ�>���:��г�iPۿ����{O�J��	�P��Eg�s��^��4�h ��5�t>��<��'5=S#H�Ȕ�@��kKTd�d6�=^6�y#�;K�3�$��C�Qm(��K������;G�7RQ<�=��'�$/�=pm����*TC� �;̏:���6�$�[�#H+�5���5�R/ݬd\F1��>iZ�075��ذ'$Ɍ	@9�ʑ��:v�F���On�x��O5�m��Jv57�e��K�h����'�.�җ��#��!��Mk ґ��L�%�v���6�SIS_-#l����n�C��7O	����H������L����"!���������u�6.<c�;�.�W��:�鯓<��u������$��h�Bh-�
�+������&�X�L�u뼻�a��c�JҴw�V�P��i
�Sv^�E��a`�S�G��M�/�ؠ2:,���c�A^�����#(�9�Ќ���%��p�|��>�A��t�e�"Lg7��:�pņ�O89}$�����l���_�o,���# ���W8m7/�t�;�� �]�vX�m��j��:�|�8K���$�tV���.S>�C�:��H�P���P�  ɟf)�,=]��������:�N�ͳ>��i�}�c9� ���:��f�Ϭ�S�@����֑���@A����t�$��A��t��Ȕ[��a��]ǘlR�cӣ㻦<m�� Gf�Z	����O�=�e�{����jR
���v�FlX#�W>b�Ht+�x�Q�h�y��J���3�e`B�9H�>6s�Hَj�e���r�`�ut����c�y�2B�C�v�Wz˰|�iU��*O��E�<�#�h�<�S�] �u�:�o�Z�.4i����ᒇ7�����;��Hv��`���/�z�t(Y�j���Ii��M�v߳q�>��;�q>/m�6E�k3����?��PCq�ngl���kT�<�-�k0��ƲG�<J��-��Ǹ��Y�vR�@�nW�_t��!}���7r&�З�N�?~r93Ev�T��� �es�S�u�[{#��л���L�D�@ BvKZ���ܘ��Z�K3�����0�_c�����wa����ߝ��>)i<�zʪB�\��Vfm��H7�ˏ��9j=n�F9������nH�	��{�qLП�8;��������R���e�׍c0��^����p�ݏ,I`Z���q,��U�>�Y�s��_$6��Dq!赁*re��4��A�0g�3��Y��4�2��˔�;��K���q���#x��=xZZZ���� ���k�� ��M|�U;Q�EF���棜9�w�^��m�bߺ�,��±h|�� +��҅'���ǿ�J)���o_MU��R���aO���\[5W<͍S�d�ꜟ��ޙ��f�ڰ�5���I!i�À�>��={���L�.0�풨��R��{cꙶ�!@>�$hl��Eȹ�Rx[q%�־�F�=L�������*�����d	A_�V�Н���]�����yC�} O`3
�s������m��K)**V/Vّ������;���Y)*b⠣�/&�C������G>�4�2�&�����}�[����p�?���G��f��{W����q��#���'�A��W��^�y|p�iM!�!�H�8iq�Nf��'��{ҸT����;V7��ʹu,K�.���q���q�#� F����*�5�"�</����I�G���I7��[BBFyy�$����@����8��x$��>�u�&/�ה�P���8�S���:�8~���4��ZOP�`[�.�Y1 #>s��=��q�ٕ�$�v!���e��i�j��Ը,U)(k��#F3H��\#:��M�����o�C��"���������L�74M:�WUU��,?6��ȳ�A��0ś�ÀrY�vlzv�{���I�p���]\����.��h]�<
�D/�Dd+T�5H��ڿ.;��? �8Ol�|9�{Q=�����n^�y�O����2-b�����ӭ��`n��.,�b���l;X��Nf��-�ŋ0O�5�Ϳ���ۊ3�<��iԔ�0A��b��ο(�D���g�Q�� �[ݚA� ڪ6��;@m����A
ѱ��hPL+�:�����P�gT^E_���"oST��$f�iϼ�>A� V��6�F���a�����jìH:>���װjG�d��!��� o��f��ONxil�z�ڱ�$�nl��jA�R�t����� �ʭ�S�����]D�3��z6�:�����S3����B�򧕈��ba�<+pR0Og�R��@�4k���z���Q��d{a��OV����~~+����`(�δ���I�`"onq�vJ�zL�U�.���w����t;���0�X�I#R8�2���(��-R����(�̳'�?�x�ʂ�2�����5BuO�'"�8
+L�����ık{BU=��g=�H���ܝ��_C�SD�6������V�ɘ���>>��sss��u�v��=+��y���zҋ8����cRW��&F���]
�dH�R}n�c}��N��%	�q�mU��k�`,C���m�7.��d�D*���W��nD�Y/w���~��TY�EJ��G7���dlR�N�æ���8��Í�[�3�������;�n�/1���_O���}$蠚��k�� �[�&U=��
ːmgf)a�.�J�Θ;E�4F�![��c(�q���<�l!�l_k����g�Z�{���ळ�܍/9���3������G�s�Ij$V�J�.�"]]�r��>+������^�(�$�*���#,ZŤ�d:���%��Z�V� �M..{�2i����9�3�5���eia��M��y��_n��sI�ːM�JF"m���V2R�=�u��;��V�9d���>�y�jo���a�;22��a��g�L��ar����E�	�wt[� g�p�[�����i��	�r¸+ʐO�K^3��s�?���<u����
�X�
E��X�HB��6'�c5��>��p-)��IȨTx?�M��~�����j-�Z�_D��"bʡ௳OR���S	�l�י�%`e�\OTYm���r�ͳ���<>X�՜E�@(!H����
W�#A3�@��w8�NcQ3��*��"1�E�g`3<<\�*M��2~x��2%з;��]�m�`��%�œ�5i�����2�%׫��q�n���U�*:e0��m4fʯ��Xx�d� ֶ}��g�|v�d>��nD�AL��q��Xa���>�����vN�	P�ؗa-�yI|~���jh�H/.�鰹e~���,̖5��@{�n7�܁���p���fc��׌ǊVC�l�;��> ��k���y,yYE���M����N{ؗ[�x�$ʏ|Ұ+�'	���X���e��eE���cϜDʾZ.{�tV�	�������P$��{\V37�|�O�DC��V�۸�h����?�o�IXH�2��ŚV�ߠ�~��J��Ψ���M��a�ɘ"����>zۻ���t��-�k�y���[�IK�Ȟ�e=ԷVÅ�����H�vx�^��?��bR�S/��{2���oWT�aT�*	px�å��:dL�t��lU���y��
�K]cĞ����{#��;��$�N#Y��pS8���n��Ӈ��]���[Y]��̑x�Q,ޡ�մ�D�z�b�<�v7����X���Zi���4��SV��v�}�����<�����@��6L��꼻��=��]���.a�=���ke��t�����gv��� �I󻱉0��v.9�}�j�U3HK��V�N�þTu�����f���� ��H��)3��*�6�N�ԆD�~'=R)�v��ӷ�T���J�^��j1舥���e\Bʦo5O���\���ܮ(X!uL�7Q�I)]���n����AЋ��9����g�.k����s��{KM]�xTB�0��sC�gk^ƎM?����Së�b��>�[��R�C�Mwc������:z2>���)��������G��\

j5�\��s�yUx�i#���ӻv
Dy�_���UHd�#�V��Q�y 9�'�Ok�����`��5kB�R� ��wqXm��GN�2��z[�rjM�5���@��[��Km���9�$V��}z9�C���ϸ�:d�S���� �^eW,\�W��#�P�mq����(cUv�V�u�!�Ѵ,tTKh��5~oO�f��,8~�p$�6�/f������Й������&J�� lL��Xlv��)8ҕ����"R_��� '���w�z���!�|,Z�MtJ���Ѭ��G��ɂ������;ӧpWY���y��{1�L3����I+�V�L?��0�~[&ӡx�Z���Qҡ�ֱ��%�]�̔�rƦ�R��R��>Ɏ�-�Q�B�K�OL_JuYT����y6�q�|����Ў�/��"<:�{z�����2r�"M@p�z����l����&B�_�	�(PO�4cJ��g�o���2���D@'o��J�I��+��xt����P��u��Й	����T�hn�P��Y̾��G�K�cb�]�C��&������ϕ<.ϱ������l$����hʌS	�8��!2���6R��L�t��Ȃ��p�g��c���͏ ��f������W�x�;��Z��B�~�B-�Lt-�xx	��_���80��<����n����e�P��F�R}N�rEFw�n���ʮ�=��nIg�v��Ԗ,�$����zV�`��]}�Z���wx)�`�����X�jf4xR҃��͞���H8�6�� *�O"�e�/Qˀ���韉7_�?+嫕�|�ج��Ӹ.�>հjo��y���:�߽���1b��"� coh�i��#\]6A�~�P;�8Գ��D�5�����.�� �k��E�֑M��t�eJ*+�"���(����$�l`�v��;��kC�NmtG�����}Y��8"�M(!h�|�7q*cI�����P�	�~�*:��Qk�O��M,�̽���y�%Te�4R�:Sww>c�c�[[�Q�K��-E���jg�р�ҡa���`b�^|�w<űꄸ��r���ڈ�˶F$��tUt���hb��/{����8��;1qJ<���7$�3��3�ե,�y��o�w-��0��!�x�h[BPT�#�=o�������$���c�]�$���~Fh����ATD�>Vp����r�00���o�g`��lޅ���3w�ξ����>Tڌ���5��(�U�x���Oe�݆%t��i�M"�3��Jv����LV9�F���'����'�棰�.��듈��� <��/��˟��?j*6���]��	򆽦~���
�2�Z��݄3=�K"SӯVJ�S9i�������?����J�����7$F�g��5�#ȫW��Ǎ��'QLљ�']�v��QAT"�\�mՠ���0u��h*l����'���g����B鬽��ZX��B��\&��6��g(.��=��)��Ȯ��VOS�S˷���X��$�̪~���aCLW8mp���`w�y�,���3���S<�$UU�@�U�����zTD�P��TۏZ��5��P6Oڼ���^��DےI��JAU��f���������nw�&��V�> Ct��c$���ʱb6�̕�%��a�@Vc���,�%��[T�����qUu���������;ڭ�s�ó�Ԭ��-�C��'�����1[��1��\�=`0�INm]���Bv2I��g�M$<��Y(�x9K����k{�2�?-H�}�t��>�BAd���A{�$�� �.�B�����fm]F�+����������J�7�-V�-E^z���s�����^�� N(�Gz>I��0>�?h����(��>9���6m4��]��)����c���ꬔ���t�����A��(H��נ�����Ύi�~�Ps��U���a8�?U�TF�C��c-�>J�I$��r�Pw�������|ut����A�m��7�d��>����W<{�ֈb�uT��.%;�&X��|�獨�E�˰h(!<\j��=h���ζR��p��E�<P ��4�o�Ѓ;��g0����M5b�PoQ��� ?��@���9$�����J��gH��Z�n�.�V�J��~���W���Z�[a��12��ʟ�i�
R��Q6��qqs�U̚VM�k��+	��⍒s;!q.�	Ff*���(Z��:��U?��'���;MZn%��'��ki�"v�|=��{b9��ϗ��^��P�B� 8)e��	�uQ�tL�	� Bs��p���=Iѐ2�P����9���"-��ő�v�L���$�M����?m,������E�R���)������u�rp�kNH@������ě����O���r�ޅ��~�7wFy%h��AA�p(3��SA��U	K���CAG��fk����t[�uGq�N�Ps����������7P���5��T>7U3�)C��(2����$hX[�Clz+�V�-�A뽴uf>�0�OZ	Sd����蘵81� J��ˏK���ng���`[���.Eh��g�*�����%�Fk������---ӥF����É�F*׺z+K���0�n\���(����zzz0���F�2*O�u�??O9M3b�5m���h'�U��v�5����H����nO�0��a�]B�!u~D]� �H�|�w]&;��n��/:�������."���S;��1�Q�-�Jʥ%�iF���$����ѬU��t�o~~��y����b�������$��>議�fV3oϏa���ݑd�,`�?�?* O�;�3c\D�j6��o����&MI���¼�FHS���l Z�
]��x�g�BMNY��� ��������-�xܹu�iߗ5���jb��+�?���҇_���}xk�fDҖ+��6Zj�;�ƻ�����ܗ�I����ii1��+��-�akkk�[.�.�:��Yk	����硙�Z��X�7Y�'نP�_u2�f7"? � י_����WN��uqҰ��4�<�ڡf�K�YTP��b��6%�V�|hr�~�E���y�D�WN��U�`XS���pne
��1[��.�������j���}�}�=���O}���'��^@vJ:����O��>�Y�?����_�X�>á"Y�A��C��`���N���å��m*|�%���X��|��n���� vu&�q�ٛ���{��ijmR߄TJA	s�B� �^��n�7!���:ƕ�h�.�D��~��,�C�k1�Vjj+ ��.R�m'���ki�+(��=�O.ua��#\rߛ�u_���/'��UCG���\�- 555:�~ϊ���+C6bgH�	�9�(�ǡn㩡��۫a���˪󵪰�kZ?dW'1��UIYI����;L�>揎�9�.��߻DZ�M�@,��S�����n� ]�F�[�����%��� �ȯ\�ĩ��'g9�Y��**Q��ZPE:���XM��a=����0����� M��H-&S�a4�,�G��[����#���A�8?�-#�7ܴ��ۥ#M�H��FQ��}m�5u�����0o��W�-�I^6ׁ��@�'O�ta�eZ��S�s�cl���p,��_Q4�����;������=��IΣ��UW2������Ux���w[�����֞�H+��X)率�/"�J)�̱���Q�n4,R_p�*�c�٦dy]{&|a� (s��1δY����S�|�qt��2�Ӛ�t ��_'�`���	�޸V,�TV��l�����:�l����Vi�q�|~}d��*����������.�@Q�+b4��t� ��3�����9�t_1k.�-���ZxçA�������0���lN،�NQ�uT�\�z&q��Sb��13�� \�ʅ��[C/o�^����K9:�N┎qJN3.�T���"e:�2���y9�$J��B��h��\��/�4��9m��n9 4�䊧���\�����L&���|(o�_g(�n�.�u���;|ϊ��_~���k�*�4/S�V�����c��t�`�A_D�;���F�I������+��/����������8�vT[�6�_��9XZZ�Ӫ���u�>�X׮^���n��9G�t�����ۙෙ��2B�������q�����O��hRNV�/����b�v-���Iޭ�Ӈ�UYIg�P'Tj�Q����n�x2�NV/:�4h��;X�ncBd3��3[Tr��2�O.�ъe;��&��к��,
�n��a���.++�X#뱴�X���U���^2����B����s�|B����7�HBl�-M;e=����9	K�����U�.g�O�����R�Fc����2��u�/쓼�]n�� @3DbF�\r�����\��Q�$)�Y��������w��^��]fXET�M%�bma���.�ToQA.g��Pi'��=�>Ѕ��zQC'绷/��DAQ^���;G}U��h ��WT��'�=��{9���>d3r$!� 8���S�o/�ee?寐C���8>���P
�����#d��Z�G#�P��$��=�HZ�u�����R����oH�3y���a��+� %U|ܾ�m�E����,�şw����䀥3)�We�g���p����u���:�<��B+�	2�c�cP�r��FDDC�&�+�Ng,b�=���p�X~�c��H����Y�i��L���Yjn�R��
�u�|���TQ�|!�s��뭴���qp�X��{I���Ѯ��,;Ls.۳�f ��?�&I^�X�6.�U���`ow��v\�C�$7���l�RKJ)���-�رEE���NAQ��y/ڪ�<���A_��C��pc�pڐ��l��ݫi&	�j�]��C�����aY���Zݬ�[8���P�]����j%��pٲ�Np�׼C�'Gz
A���{I��an����lʌ��Fqm`���7���r���Sl>k����x�[�]�q�)"{��t|��O�%<4 ��I����&aި��� ;y���=�z����r�x#�2L(?;;���7�0���vv~sE�7R�r���r�D�����!�_<A�>Ln0�ނ��H�-%{S�N£�/f��Z��q�ܤh��e�����ĹҖ��]�4o����#����D��N0��u������i|7��.�A�
Ң"�e�EW�������o���Q[����OY��Х�_�)W�r���w�3���P��g��?,ɾ?yһ?�&�����_z�B1�[7�<Ҧ>aǙ*�N)��Y���5ܯ���ߊ��R�]� >�p����v42��-����
�h����f΄
E�1���h�� 	mQ�A�� ��Uj[�xdI��|4���o�63�|d�[] �(���j����]�f��[α��$c��X�o�6	8�]�g���F������2p���q�pFnR��r���PT��P��n�I@�p-�p���x��IyE�vw4����'	)���SU I�̱+uQ{��W�U�RC��`e�v�OvU�&�np��e!��i䆺/J�Hӻ��(�j,g�K$ι�g�"��������=�85,��`y���Jp��`�������� pdS���]C�jR�׼Y$l	{�#�c�T��!J�]+��g�%D"	�"��(��N��
��(&�Zs�q��C��aA�1UUU�9��ZN�$H�=.��%f��R�m�4��!��ᴬ*?��@�]JwQ������M\�<��$ѯ�1^�4b�أr8b�#�]���ė�W�ڭ��G+S<K�� �Y�#Ē	���9�\�����@�$���G����'6����Z������-���G��a^�����bY*:]"����&-�H)���%���e,=&_R����?�9�S�����ZP����c���&�!eTD�<`���$iE�Y��b^8^���օ���^�۴�b� ������L�����ע��.`�����E�>�M��i�m1�1�;^�/`ZG%1�m[;Ch!2o/����s;}$�W��ȩ����E(��E�z��Z�YI&����`^�7,΍.�G}Bn}CT��S�z`���^ 2 _���[n1��&����)�.�U��HFy4j ���xT}}r?3���$�y���f� �0��L��]tp�A��r�R(,z��U@Y�*�ń�sK�!�����vg�`���y����jF2ݬ��K݊��>bi���g9�i�r���Ү�p�M��|(��tΣT>kz]�\�G���N"� K:�zr�r{i�}�����t,u=#��勏]���,���"�we�����'r-��_��8���c��@Uֳ����
T���ț��?�C"+[J�G}z?�ك���/��%��}�bbjj4A�Y���*��|8c��A��໬�[j5�!A1�&���̯s�x�8Dc��i�����YTf�4h]�h����I������&�B0y�KHlP��"I���4���I�á�֢�!���v�n��v��jY�)�b�Ɯn�?�������qZ�⯾��6,�(�M�}-3�^;. �T�쇑��b~�M�v��O=���������-bf ��IMH�������<P�
����!�Q��=����Y^N�~���/�t��k�.���*�=����z?sIg��B�:���e��ђ�Z��?DQiow<������Z�X����K���?��%�G�˟X�wg+��r���(�L�ٙd�-m��2n��e���x�և�[^4D�l���b(ُ�N��6��VoH����}��W�����Ϡᤚ!G"�4D!�룬��� 66̢R�����d��8�XC�Z�~�NG#��`Zߞm�u���W���E3����[��8{˨���m�Ѝt	H��J#)��tww���$���C7Jw�7��������8á;V̸�Zך�χ�� Z`80v���Gō�r=^$�
�㤟����_��EE��(zMP��(hoE�咷��Z�vs��a�-6H��:C
K&��)�	k�aLA���_��<vDͯ���p�]5ٹaD,�+�#�����6�D����Sr2��O\<��9���F�>`_5��6�@�a�����\�_�2M2�:�?.�h��ٜX%;w��Bc��Gc�/�v�K5+�@�* �����n�K-����uK�b �>�;�j���2_J�痃R]��4���2Kz����x�U���98<S��d�HL�6�����S����B\����\hd?�#�'6�1#KI��(����Zt7|�<��O�$���P�� ��m���n��_2K � �S�? �0!c��P
y�Wf�������>�בN;�X�)�-|�$S�er��~��[g�K�_�O�Ȉ��>���ðy����H��_pI#k(���Q���'2�����V�;��ľ9��,mH
�����P�D�`������_2Of�>��tr2�����P���ӛ�,�� ������M���)���>���/��:62�(��+$6������=�o=|pl��BB�]��v����oz
K2�L_��dS*�q�p���D��~ʌvL��eZ�z�����J�DcJ��Qv���s���4��0%�%~x���!�����Nb_2~Z�B�Qe!9LA�������%��̩8�=�㰲�
B��h�.��D3�ʁ���b��D(�ã��X>J0z��ۨ�4��]�߶���D�85��|v�����x+�RyQ�}���0��L�)S�~x$Q�X�3��{��ʇ�����B%A!Q�ݳ��}�e�K���������L�%���ibE������l$�./[pv�3k����g�����5:-�p��P�a�ŵ��2�y�����36.�'�F�˜�$��.�Jm�m:�(j�����B���P�OL�a*,)�,��c�c��dWb��D$Dj�H2y�'y]��O�����Ll�̴"��֤��c�M�3d����8���8�a��ي�D��l���iX&���Q+�=���ؖ4���s9�o�5�L�8�^�bc�T8��~ۗ�J~1�8rZ�C�d��TO綒���UJ��Ǖ	z8�!��Ƃ���Y��Dz�9�~(�h�q����X��?�t��s�L���s��Xv]�݌eg!B����]�E�"����hh���J�2QT�L�9��,����Z�M�'�9t��0�Ea�"��J|�G��������M�S��7�CS���ӷo���z��y��:5�o�m[9Z#S�/U(\\�kY�������Bɓ���qb[BY�����y�z1�Y^qF�Ǧ�`���g^B7���B^����9��p;y>�.=�\�U�	�0��F��y���+���Z��i8*V>Ѿ��e��i�ީm"�$K/7X��k,&����X�^3��oڥm��� 3�$Yq�a��畓�ñ��Z/��H�Fh���hP�܆+���������6D0�Ba�e˛�:4&������Gݪe�444jۮ�5�"�5��L/�[-�~*�wl��^���I�/` 6|�T�x��!$q�
I}���ψ�P-������*��GEB�����{��Da��r:��qn�<E8��Z9.W:�'��E����u42���:�Wo�op�yuo�������N.IRR���MM'����:�=��ё�A����	�I��^�X��|"ݗ��i����������ZW���:W�'�kBoN6�
�]���[Vͱ����)>�Y
�u��X��kb6+�a���zQkl�y�������S��|�q�o>���U�Cт���N6hֶ�vi���oQ�R��Nq�S�]�]Z�
M��Z��Ĥ��rH�a�e� DUC#��"k��֖���@W=�ne�0��ð}&�^\F&�\�xS ��?C%V�e̶qbU�Fxxx"��Έ�}hnN< ����Q�no�hh���:�hm1���������Tg}K��?���{�me}u��gqe�Z~\�kW`@_��?KD*��[:K4��u�����ܠ����	I�.H�P<u2��c���:]*7�)�Q ��GKO�x*je�1<�����':���Yt��
��+!�a�����ɠp������l��>aY���&	�+���܌�T�=q����'F��.M~zL��~.�8�ʻ��R�<T`$/����KJR����iY�=�
<�l� !�'[0!V<չ�;)QHim��W`��H�# ��D*��Jq�(g��):�B�|������������nj�E�E8$!		8D;�郛A��k�V��v\\��vP����c8���pU5j*΄P/�`� �����O���Uvyz 5v�xw��0�.�c28(����xK�K�n���ۣ�N]DK.2˚�W������P��չg(���4��V�	�Ys���c�t�t���a�#$G��fp|Z�o�'2����!u�7;��,�%�$�ȈH(]���9U>�Wu ��Ǻe��W�q���R��=_��	�� 5��Ρ��� ���0ܨ��t�b��t�N�����yҰ�?��b������ć杀������ף`�~���<�s!��u�[��9\ZN�>��E<��N�{؉tF����޺� �g
E�?�x^_כt�0�I`��Z�6���8Ǹd� �=�˖�5'*2���{hӽ��_^�C���ٻ�k@��Q�M{��_N�k����	4������Po����I7���?U
���r�{Ժ��S#]+�mjj�OG5$(^�59zX�q�P���J�dh��[�Rh�������������O���Ս���""���[pc�(Q+�3��E%�:�h��6�'ґ�{DFF�D�Uk�^܇vm:�G ��:8�l��΁���u���J|���Jme@ۚ��g�!�C�ULKq�f��-t�|^gLsu�y1�4b`��{�,30�;�FDaJIxP��r�d����f�K~}�Q��g�ħc�ѿ`��:}E�MsB��xp-�}'������&��`ϛ��O�;���vuO~��0�ګYR��m@��qr��A�o���2T^r�컢�2����+%a*���I�:�[3j�(
omM�ȧWX;����d�OĦƵ�V�[-s@�C��h�e���c�)b�)��{�T7�3�D;mY
+�%��o=� jnOh�׾��{�)zY�e�a]}��Hn?"���z��>�@���Pv��]��d�T�Qx���j��2'����t(��ɭ�e���ɱ8	�0*���$����5,-U���X�"�;~U�.'�DCÊ��W��;���@I]?o0�?�vj�7����tJ`K&\��j,-�<�j�6jS�4K��.�`Dkd��9L'B��;s��lYT`�d�q�7~h~�9y����Ւ80�K"P��k��@d��}�Ϲ�`��2�#�9�O}�������/�;B�a_�045��mP������L���
����?��#�jf�E�,p���e�]#N�an���T߶�ç��Fu� !�[m�����Vt�eQ:͇Y����"�@E=4�5zF#h�m��)�����ڿ���]'��'yQs/�Ài"]@Uf�U�0�ƣy&���±�<9EQ�?e�BCCedd���$����o�̧�ڷ];�]so�a�b�_̭��e487��
�Ṽ|��Yv��Fv`\�_2Z/����E�Od3��l^0b6�¿�!*驿���^��H�烬Sg�d���}%RcGvw�j��	Ab�R>a\�RO���R��g��!W�T���]�Z�Ơ�Be�m��°/e�x���A��U���K���f��.]~љ�p�����ݨ�ە�b����P��?(�����DP �ZL*k�*���RF�|�co�>�����ƪF{�c=�B�t��)�ߥ75cV���0��ڷ\��=��k=�-	�ъmH�m��ͫH�/�����}2Е��O���GF�`�c��1��5�M5�l\mD���أ�Co��}��^���ڽ:x8o�L��_����f���Ylr��:�5��߳8�B1/}+�t*����1Z�U��������qf�-|3�%srs��;p�.":����u���֖�����wo/!��� C��ڞ���-tg<�,y��+����X��i��������_���̠@|�yrӠ�V��m��oمvx��!_���]���\�]u����wP;v�E��7�K>_E% ?b�?WS1��%5�,c~-��/��i>п�LNDA�����Y�r��>|`F��.�Q�$0ƽ�/R���f��) �[v-M�&ZvM�
L����sV��`B�0��*����h��Ca�35�?�'��H��y���s�! �-|k�rX�����g
�^���DW?��t����e��g  �
f+�c��T& �����:1��nH�+#�s�ϗW�ۮ`�J��
#c����ýf�3�������[�&�gXX����-��`*l����%�𽅒���+++o-����"f������]p����wo����҂��CH��z�V���|F��ߑ���>�bb~�G8;�k¡�] ?+���6�/��2�߅n*�럞�.S	
��kO����,g�޽�ĨAr�k+tC���<��Vp��/�}���&I����7<n#'��n޻��S2�F���!�����t�{ק�a�v(:B��i!�@�	S����pz���U�|���I��p�b�tss�tOo�>T�����_s�D�}�6���t��O�*{�/e�nX����|��I%����)$��/��^-y
�B?���Q���<ǃ�,�/����	?��������	?\�̮[r� X��x�l�(��%R!øY�^���ܬ�h�����*�c�*t�*�j�Pj;�|�ϗL�D�{�o��ZO�0���3�Mv���'�e�q%�;��o��!�q��t��Q���M�{�ܹ���X���s�.G$n/G�������Y�:�'�Q�e�9��gJ���V��3�*-�Gp|\�:~����n�k��GhA�����@�#`$^����n�)r����6>+�O�tZ�<1;�Ku�m�Y�F*T�	������P��5=�vmL�'� �ŏ6�f2��uX�窆pmM.�����yIE��o@���z�; �v5J�֬�%�,���#>��[��ͩ�Nۄ"<i`
{������I�������_71���EE�3)�vwU#��0Onݡ=�P�	��3��?�ak!!�5�,\�J�����`�y�X)�j^.y?L���k�#5���]�����/˿��h�ϟ�ri�����L�-X�5W��ľ��w��܍Y�&��Dr����0�x�N���a�Y�~�����~��L�͞��>W��xGv��W�HϾ~%ADB�~�jiw`p"&&F������]���e������o���XB}�y?~p��n��O�� <�� I��aL����:�V���f:��D�n'nd�c���0���j�R\Z)�ܱY�mO(�m��u!����<�g0NK�����o^���pS��s�V�u������%B2�Q��a'�@;�N�h[�*OJ���[���cZ��d��hrC�O�Z|3�4η�|n����<�-թ�y�f͞.�
�]�@(�(O�����V;h���䆍�$ "��)��5�����6��Cv�J����k�ī r�	r]�wԦ�Ub���N6�E��������$�Ov;3�Eq�Ծ����YhPۯ�ʂ��V�!
&%84TqN*7d����^�����������>�O�������R	���,�?�j�q�������T��yJc�h�߽���!�]:��_y���0??)��RJ,���������mi�5�~�[Ӟ�ݝ����TH�A�s���e��X�S��A���������}�7\`/pk^�\�O )?8�$N�ӭ��Į��B���_���Ha��GMq����#y���ګ�f0�P�X�ba�����qm�ʴ�C7X��� �\_�=�:O����?��)O9�������"��{?�J�Pjw'P����v,t��^v�C����\
��+Ć��mN~��M,�֠dL1��S�(C�7��Wp�ެu(p��X��6�.��6JT|plx�]���ۋ���mj}KK���28��-\vFj��!Y�¾"�톖��!/�n�
���{��	G��� i�Q�,f�D�j��Z��%%��� r\ߛm\� |��L%���Nu!�H��	S I��E_��Ѫ�)�?��W����1�9��p�Ui;����v��!@�$%�C��*sj�Y,������ɳ(����PU� b���o+[�BT����.��G�a�^��߭� YO�v$���+��+d`pT�a����檥Dl��$�Wo�>���{\��Y#���.���m�r��ew>�e���\����{������l��P��iýb3iՆ{�a��@��*��P���)"����@���1|w��������̀��1Ǥ�9;;\~1��L7kStV8����ξ�b�7���٦,�c�c
xOv|����1��%�F��ǀ����� �A��{��i�J��[)��
��m�3�vM���w��#�F����5jo
�+��iI2ܗ"�@,�lg��:X���
�u�-�Z+�����z(S5�񴺁e
u:a;޼D;���N�1�3��;5gF���m)l������͑Kֿ���\W����:<���JR��x<���������v�O�Kd_:�TҌ?b�iyڨ��ɋ�l��>��/�H(����z~�#�i=g͢{�#dH�	Tӄ����N�����W����6!)����qF���Nv]80LO�X��J��\(���_fX��JͫW��y�g"w+N���ٗ-.t���o7�֜�8��.�(wT=��rq]+��A>��h"_�U�kW�br�X'�@fR�T��,�a:��
�ˋ��m��z���X�x(T�c��:��u>\�[ы|�rr���Ɉ��}Y��H[�����l� ��f�a�޹�����U�O��8AP��5o�G�&/�0��Sm�˵��>�9�U�x��V�_(��_�ڨ��������`�\�~a��Ô��Ht�4���%�� R���j�	'9����*d����.Ո�e|�'D��ϒj��w�l�(�k��{��P#K�ņcR&+�p&�";LiW�@
�Cr]��!��0�	A/N |���z�������� ����-��;�2�I>	-�7)�����a�T+�V������Fe�Ve�|����Yp/��c��j�:�?d?sz�Y8�x���%w%��:8�_�R���w�4w��~\%�CF6;RY������������7��2�0L�����f'��v�/��"�����>�ٔ5 ��I
_zqr����Y��	x��X��pG�����__��&���3C$��'=���A��5��ȟ�RB��T�x��%I�"QQA�\��%��@�H�]J�����#�&��(P��v�agǮ2�̗O3u�oK��}ys޵�LȨ��cм����(�0���x:VE��u�>�/���W+�OUx��ݜM�c�B����џ��Tn�I�P����^���O<����?�p���3Hcs�޸S>��*�m��9�����5 �`����+����}��u��̸/������G�)��~�®[J`��_(enWG�g����K�B�G���H�R�D��V�I�V��U�	��NU���µ����Th��}�Hb����
����A����ao�����zjj���:�}*x4��$���;�@|�7�l��b^�\���i���	VY�.!����񶜮�hUkr�Y/�g@RrHpW�����W���diwH~���,��C��,�����D��ܿ���<j�	�[w�_o��N
�� �@��ɘH���K������#���/	��YX��o$�D4^�LϿ����S���q\>�Hsu�U�H`�K��[��ˈ���!������HH�����q̑��<�������U����F�ꮜZ�? ��y_�ɕ�S.VL���S����2���t��tK_ֹ���~yE���P������:�qْ;M�Z�ؔ�+�<�g�����v�vU<*Nc,.��,�ێ*jP 0!ecݞ�τ� `"�s�A<������#��;��d�M&k�#���>�e���AV�~�%8j��K/�.�(���8B0�k��CN�BF�����.;�w^!�Й���A�l��~��oYv�|i�zfP)�HqCw���NK�1 �V�;���4�e�g�+���taA���;,�w�2s�j`���N�c�[���9�y;��T5��eng��ThM_^��]��JŴH��n�G�8�U^4OZ�,eg����˾_�]�������msɽKW�}����a<��	�� �t"�@D 𗏧R�k���eL��ھ�Ϭ���jx��I�و�U"7�[��w~�}./�s�ǚ1?�z�~��K�t(�'���߿~�M�0��elbB��y�]�eX7n��j���~��on7�#	*�B'Q�3�I]Q�N���E�l�uj���˂^��"�W!t�E��*��C��2��Ϭ�O�Ջ	===#"#?��1#���>w��r
		)�U�Nܸhb� HmX��U�?��_�|g���߾�*v5��!�v��^'��{�CM_?�]��~R�[��@F������|hӯ|���7AĨ����G��O�*yh_��8�s���8'�ϼ��?�ڥꐣz�yg^BEEB�Jf�;�������&��?�D�ɞ�ln��Byx�{��!s��?���(�?C$kw��
!G��rrr���aW
�ա�r6	���4�]6`���`A���������4��R�����]�X]%���k:z���ϟG��ͭyb��7�r�j�4�d��Y3D������/����W�IV��¬�m�MDl����.0�/��� u�2�2���F.*�ɣ�33�q���o!�����M�i������ģ֛��m�eM� t/��̀x�>o��B����dՔ�g��s��'�Kp�m2�����թ����)ŭ|qUB��ZVÎ��ir��6���A|O���x�֔G{
l�a����������TX��5>gk�^�$�GIn,v+�׫�/p()�Z���\,������2af\dNC�0��������t�D��Y���Z�a�;##��u�a�]���D�?�]����@��Շ���B�k3w:��*�S&M�x<�A9U��LJ��9� �_��ѣ	J�9n���\���%���}��{��r�i��R�<�#"��s�VW�o�LL�O�:�S�b�c_AZ?�����j��jc�[	�x|��9�&�N&�N�Ls��R�h��w��y�6��
ǨϞ��
��ǂ��ǻ"N�]�0��,O�jmI�{�Nc��
wJ��yK�	d��iQ�h�2K��	��Sp?a�z[_�J�m�=�Kb�P4�d�hZB>H��$i�vi�$��[JH������E�QlX�'H�T�ʧ�ɖ�t@׺ϟ�n�,⋣B�@�P]�,>����"�þ����l��ˡ	6[� Y���1ڮ�u�3oj!��L���yu��
��jW��J�!B	������ppp���0)ߒ,6��n�~R�����)᭝���v��Z1�c����ؼ,D�-���G:�^t�d��\8�ԬQ
.�97(o���Y\�_X��@��P�8�ፔ�̣��vM��p>%��'��s&�A��I�k�/O@�o*.+��=ocnG�3H'& X9�K���|�z����v�+�N� ?���ts�����Ϧ���.�������,_�`�`P<��.������O��@GF���99$x?
����[׉2��Q?���S����Uz�Ƹ5�;V��ڛ!�M�c��	���})��VҦ��÷ �Ѽy�_���2��] 3m�"���/y�PSS_]�=.����K�},I2M�!�W�R�=	�A.�/�>�i[�b>딼��{��@A�R�5����G����C�x �[�Y�� ����GIA # �h6��466����&
�v��7�^[�ļ�v�@�ft�w���'���'�fW��6V�,��5�׬�"�؈?���֑�%�k�����Aȉ5tb7m�K?b�_�?7�gJJ�C�U��;������h��no���&� �|��^t�}��hV«����������`AK6�����
v���T��]w�}�`�{�z{�\.�X�`v�����g�E�������"�����Bܰ��T���o�!�c|Ճ ��f��>����ҷJLMaW���8�۳�wL,,]g����<�J� �
��2����A�>X�,�Dw���G��MM�G���k��M�K�Sv���r�n�"�%x�%
�P�q圦��g�h�7Sm�(����7o��6�x'�_��h�0��ND�z�18���*��|����y�H;���G�FJJ��6�[A/Ь�o`r͇RCA�G!��/�.�8��2���!�������؏���RU��_�3ŗ�9��+�(�X��oS�]Dx$��G�E%�C��K��,w�bg	���Rm������ݗN&�U^�^�
���7m�J:G)��V��+�K+�X������43��Y��:X����3���;�Qq�"`�#"P	����J[�^�?^���Ef��5H�t`���铹fb��*zZ�T�O'��Lrn��- �Nĭu'��}��w_�f�ʶE�<�ؤRA�,=��@H+uji��&o57^�ă<�+P2����r��/��D�٣r���j(����aDߦ��(Pe�k���yߌ{�:���֑PS@8����f}ᡂi]Om���y��چ�b0^
9�����u��X`w�l�D�[6ل%$C%����Α�_���ddP�v� ������E�	th��0��2:�eRҗ�P_[uKII�2̿��BP�m�\�
�r�ǐ���&��I��]�ŜI�a�)T�S�S�����X�<���	����p�^xD�]t<�N}%���49yV���W�PA���`�fYl��t�!�VS����~��hjf�OY^_Or}}�T ���	
>b�w�{���牉��,Fx�W����3��x��ȉ���.��+'���/|��5����^�v1F�-��H��ÑB�r������m:�ī����
��co]�
�53�����d�v��ز����c[�ca�V���m�ُTn�M��j5X"�6w�'		.fz��9N�߿�%"��,����<�C!HĢQvv� `Aã���_f��y����g[D�	��^�p_��%p+���ȉ��Ad�E�	����"h{ћ���X|v�F$�a�e��v�P�Pߤ�(����O!�XW��f]ĕh����+n��QB�Mf��QYqc��`m'e�P7�e��������"�w�Uݲ_���ܟT����.��C��{w���G��S3:�����,|APW���.��'�g+ �����{��7�8��U
��U�Ht��R�w�F�;Ώn%�(�>�b��h�p2�j�Ң"f��cůq..@�$�e��F����c��=������F�.�-Yp�]�R�<��oW���|n6�U���wğ��+}��p��z������x�2^npp0xb[�/M�)� �Ԃ���b��N���p9�s��`�����vG811q�E���
��{�Ɨ���b��WӺݲ'yx܀H�b���* Q�XO�emD�v���ȩ�z+@X(b�oF����>T�WU�+�Q��u�8G���R˯�����|d��R%s��! ��9�v$���_.�٩���P11%tuɑ�QƀU���H�M��=�p���V^�֙�B�&^����E�b��F�I�<��c�[g"��B�n�\�n�O�M��,*Q��ځ���76LɅ����#��]����_=�su��Z�|�~7V`��|�v�����&���ڊ�8�eZ��Oĕ���e~=�DBB��T���mjk�+�n����#?�mhhĝ�mӂK��%W����}��C樱*ELNH�FyX������1��pva�)ܭ�H^�?~Ё���]ZZee���5㽹���R���zCG�Xa׏���Qv�zy����:��˰�����S�H���B��Fw��|c;�f�cc|�=HM�/��
`��^�	t_	���vΫp����n|F��hd!����{�.J���q�/E��E�G���K�D>rv��kl��o���z�C�h]
���L
�?9�Rp�{��l�q���m�/�l9|(�J���8~��(�c��ڵM.�Ι�K7:t���5(�O�Ku�}dի$ W�B���QX�	_���Z�Pͪ��S��Ϛ���w�;"���*�ܔ��,?�8Ŷ/��������ƚu�S�I2��q�\�}�"
=+g�g�<ɐ[����|32У�\-��P_~�Y�����U���3XQ���  ����^Muze}�_,%��q��%�3,%_L��t������㰟8O��׳�>/���A��p\���j'�ڻ߻b�}�ƌx�w�LhҍF.�3��	cTB�-�}���
�D��]I�F���Z��On����O�x2ٿ`̪w,���A�]��� �,<�Ŧ����
M�di��{v�p1kO,�{S�F���D�7��;��b�ņ�lg�2r��
5��ʧ�����[ݗG��:ʯ]{��m&��PG@+�V�'��<O+�,�i�����[ɫ����Oj�x���6e���W�hj�"�`�4��}I��>5r?� �����L�����@&75�i)�캚y��~!߾Q49�Pab+>��{(��^��Ь<��j{Ϗ�L�:�Qvx�U��TqM�9�>�	�;/	xFB��@!��m�c㿥�Ҵ����+LF�$�A����GK���#ɚ	.E$��0��T���y�TJkE�$ԡԿ~a��1DќyaazQ`z�q�����6�<ϊ�o�yW��v$�EwrV�x�D��-_N�8)eD�UbZ�����w�ͪk�Ȕ2���؎�e����� �4��"��G�@$/�'�P��	�ϧ��i�t���_�!WU�΍�������Cd��@!`����!aa��<�v��@��JU܈�������
eș丟^�|� ��*�T��r�`�6�b*8x�p�h�����}�s6����&��E?޶=�L�D�v�Y���d����n�Phh���	�״O/��Il��,���w?]~H�n���OĪ�M!�m�g	+���� K�ʊ�Zo�maY����c`pPY[;J�@�ZD�M�	����ivs�b��$���>Ut��7�6e-�ecfF>80�x����ԢSSq���p+))A�fcZ�/��Ջ%--�0�b�h����o7��Ҋۮ��U���P���!��)�Љ��gM��
0�V �TW�6+GAB�0}�1R~�!*
9�^(Q�5�n=pn0�)�z؛��Xe%&�+D���|zz�V��1 �Q���|QD*��F�M�Ԕ��h����D�Q�ls��DDll蘥�@�X0|+�}��6A"���ee��M܆wױ�~c9�|�[	�*֯A2/W���Ā(��ֶVZ�d��y����7�,6:������[.0Z��KFc����?��45�Q��J�u�F&�_�h���߽��b's���$b�hLF!!#� �UA��l����q�~�y�f w�
U	��.x���@��@��С���A]��Q�'�_����F"Y��8����R=�T�x�Swjj�V�@?��;�x��)%����l e-�,��X9Y�����&K]';:'�Myk�y?��taEH*[*}�G���;�?�	]��O���DW��&�� !��rR�"2�(55:`�p	Ic�"���	����G	:�Y_�F��(��9S���e���ĳ�Ѷ��(;Ĥ�֬%p#�?���������d���G�+���z5NOpvҔ��:���F���{YM�j�5�B���N��A�\�x��A ����76DI�NZ
wA��{��c��in2,`v�n�X88�%C�}�-�u�'��Fh̶p��Y9?��E����^�x}q z���Z��N�`3�R��`�/**�Ɉ�������ʯL �f�|i��჈� B7grY�� �4	�ݛq����>G�	��"���:Zzz$�R���f�ӣ�ǻ�u�������2Wh?��C��\�\�cA��5�u�~Aw�_���!���;O��0��7Oc����ʞ ��	�B�F�S�Aәf/(a))���z��
����z�Ty�6 �ͪ�H���ִ��=�����&?=#����2"2'���g�ց��[�3Z̆��}Pg1�jg'��=O��I+!lkw���7v	��_��4��I\����w!�h�;��Q�"=`~���P*$&XL��Ml ۾�!�D;��r����8�K�Wc0&����ɏ�HJ�ֶ�m��`��Ľ|��[�(,F�L^�8��Q�lg�|V��0�t���y���w~F=׋�~� Va)`PCgm/��>�e��aݒ�Mn9��srs+W;��G�9�Xyc���b}��.U�7~h��	��>��a��[٤:�ԕhk'��?n5�H�2���l�9�!����{�644b�a���=Y#WR�f��7Z�w�\v�
�"9��,k'HY�]�-�.4q����xV��i�2�|����40����g�y%j���8\�z ?����L�jg� hD�H�VӻJ�����Р x5c/�����8�`:Y��Lqy+zA���ż��r��q'��Yc��i
�$�I����y���I >�-/<lD�eƙ��<���5�v�41�T�Vdǽ  s�]wǉ.Ȣ.Ef�v�7�6�����h.�fsš'}�O�$ޞ�y㱙��	�����?����`񹬬�f�t��\1��a���4�V������;̪�ע���!��Ov]��Mk6��tBmk��sZ���W�n͆�/�,����'��vbDI�Λrw����3�&Ǡ�1*����JW�spyI(�m'�����d��]���|C}e���m�&4y�?��NS�ѿx
}�N|���prJ�.�ʹ�S̿{{�?i�Ɛ�a!�r�����"���U�S�)W���?�]�,���l���1�����A�.�/�5����+��.ʺ� %��mG�������_�𗌻s��}��ЏbX��5�v��E`^.�<�/zڝ����'n�CG�lֿ�!9��N0;S���/�Ĳ`:��vѤ*r5tW��j��y������)�,��k5��bR<�����<-
т��R����YS���<?WL����Ia����j�y%�q�_������,墹V7^j�) ��ΜF��OŒA}䶙.NcG��{��rj��ţ�Q�cjP���KE�Hp�%��s��\pp^�eY�/���<d�ո�h]��,�"��V�L7�#���{�W�TtwP/�7&���Մ,��� n,�}���-�]���n.�)w@���Q,a��N�rL��3�--�Ǿm݃�����>�#=b��A��wҙ_���=FE��rT�SbB���� ��I57��y�#��[@�^l��"����Q�30�Ag�X�S~3�J*��\520��z������VM+�! �L����+$V*8=�\�������'�������O��@��,º�s-_�K8��T���Ç��=9Yp�'��G��yKl����H~����GlӞ�#Tj)� 6�_(�eɨQ���D7�����L�[(��Lz�\'�=�Ƥ�2Z4||$�������i<����(U#O<�D��`�y&{��#SI��G�#WK�ՁH|�����g����*��.�)�����#���w B��z��M��z���擏:�\��ɧ&�_��K��~�%�y�����߮��p�ֽ킇�/���@�X�M|��
��F�����>%�v��z�_��p.!!RG0��3cA�v6L�y5_1��IJ&�׋���?^H�B���U2���!��f#չ^��L-s����h�c±i��P�rz�:�Y�˫�@7	ˈF�f$�yD�*J9�e6ޞ�j�"��Dgh��ww9�w8���H�@6��3����n�|@s���s��>����$�A"S�q-M�}3>nQ��n`	�M�*Cs���J�}�����z���]�-f��$?>Y+�y�|�����:�J��6���x��E�n�~}SΒ8����u�i��rv�/ݤ�Bu�*���7�CW2�)�|��`g�1tb�h�IC�]��53&������3��eT�D�z=��H#����=�#W�ZTJ��xD�y�O�P���h��� �Ph���7�il	5ը�~pD\-#�¨+�-�~��N:�K�TIa �����	�j'O~E�F<1��f=zB{����j�埄Grળ!~�'�:E�J�HeK|��8�\1WW.<||�K���UL�*^��񤃸L��o�Ԃ�ǫ��0�e�p���.W����/��%&�����IҼeU�U�v�?��.Ux-��q6<:5�������OҔY~Q%%�w'�3͞o@�Y0�3���P _�Hcm�_"y�z�ͅ����{��T��G���+{�5v�����Y�_a��x*�)))u�Su�-_�P�>W�&�r�L�u�
�1=D�[������<1���oF�"R&�Ix�ɗ|N��4�[3��rHm��3���KQ�Szj�2�N8����HQ�u;}{Z�������,d���P����z�Ү�s�B�>���|�+�r�(��Fˎ���zE���=Q10�V���� ��ncM���y w���]��������YcM���G����U@E�>��PBDZJR�CJ�AB�[:�K@��A�n��f	��������Y�v��;��33��l����ᴞ#���]i������t�n�����5P=//7]�X�/Xi�G/%�:�ܠ�+7��,�]��`+�G>�ogG%.!!H�����Y�h�Jē�1�.M�CB��n<&���Dz�:]�8++XJ�d��
&T��������v'����=Ne���!3��R��+��+pct�)�.��z^���"��@t�%J�h<�3��/��'��B�O� ٜi*5Z�|����.���m�����{�ޣ-��
0��D��{VNNN�P�y��(n�W���~�>ujN�=o"�Ng�`E3[�:]Y��t:&S>��ܔIvj0�o��6lf�����7ӈ�����D�����z���E(�4�7%��&C3����9�^RsIX��"
�a�r�Z�k��R�U�'���a��i�״L#T!c������lSo��SQ3�^V�f��Քϧ:�9�IC���lZ��{g�bD�<m��>w{���������T;c��_�e2��ȥ���3�����;>�9Y�pn
����Z�O(ک0�@�yGy���y�Zv*�:�q�Q������Tİ���
|=�L��������-��u�Ty�IQ�z�#M�)x;rB�߲��m[B�m� <]���:n!T�3�����i�X`��,��4ч'x~pOrn-���5�#
BVxM�&�|���-j~��t>�N�J�.5u�m=������J��SU#����Z0�s�bO��Ib���S5�Ǡ�b�� �ȭ|��
��P���o���-}C?~�4��261���������%Н����F2L�:��~���\�;n�J�|�h��+�V@&����NQ؏��y)�F�:���*#�}�/s��P1�?L��
����;W��dq��������íϷ��LSd�K�.��^��E,�q30��t�U}�j
���+���r<��b��"+	1(�����F��u��� Ǳ�p�9�3�������s��oW���"�tU�\A��eb��+�8�z��:-Y�O�B�R�TW⊘�����������#�h|�a�w�M�7����E�+)��گǤ���{�a�������)M�`�p�T����m���X�N�I:K�يě����L�ܣ����Q�A���>������߲��oA��q* :���+T4�$������Q�UC�/�-��-#b��?n���_��o�־�0�r�@��(���ѩ��a�}�/}����׍��(r'����M�飢�g����ZXX��ٗ�e���ul�Iw�Z4�o>��D Vʥ����s�%_�N�L�4���~�r��@�,V3,�^�<��Krz%O.� �Z_���g��4��V��H��;�=�
�����tvm-������5H�
� AsP������:��i*jjC�;A��予m���C�� I��P?|[�m�� L�M�>�w�yJ&@��F^LM���Y�w]3�m&9�v
�Sk����eS-�������A,��Voo����0�	����}��K�D�W��s�/�#@v�
{1tI����o= }pt����`����^��0��(��C��j�������^6E���-�%FGF���V�-̓��{I��($�а˚�4�e�����t�P����.
�H��z�8
��`�M�fY���Dn����־�u���z�Qoh�n���V��?{w�u����Y>�ƙ��)�w�gp[��~f#��u�ݹ��Ъ�N0Ix�my�E��;Y��LM}���5]������D�t;"�sn�]��*,"8�Xdd�33b���o�>wi$�F �ՊqM���+������ ށWdd$p�ll��o ~����e倹9����Zs����ԯ��(89񎏏C���K*�ٱ��" @������J�U����窱�"E�&)9YQ]=����E��䤰���_�`<&$w �Yq&��F�Z���v[� },���q�����|cCޙVQQZݢ���C@^���ﺽ:�s�'$��8���!y� 6Q8�Ш4F�?|�W�q���f3hKy�(�ZMI�p�&&'�W�ȩ���<Zn����O�媻�C�e�o�p��a���w1z�?P������U_�E���J��8� ?��� ��]<�N�N�Ȉ��7V�����,-٦/	 ����^j�7M�+���PN��blן��yf�������nuAѮkU�x��=�H��B(3m�w6�]q�����F������;_[_�����v>���jx{5S�)��d�C����XФ�,p��p���|l�z&�Բm`W�p斗`A���ʪ�p
�R�P}�P����qd�'Ы�nn���&��J_L�r���:h�f�� 
E�HB���L�(����{��;�"��;��\ xiii����
:ߦҿzձ��MDd�Fѝ_TPh-!���Ed��v��W�E'$�j���8W����F%���^��Q��/&݆6�:��@nn�F�w�O��m���@"�" ����(ɜ��s��o�k��U]z�7p#^�q��5���uqEi���j��ј���LOk5�h�d�,V�ehl�~��c�L̠��NE<wr͉��]˾���=�G�V>����)L�E�3k�����y�����L3�|n������R��ő@"��V�x����ʆF�b����D��[n�F����"MG~t��W�2�o
���s��_5c����ȃ�vH�ט�%v�F�Ɉn+�,*�Zj��� ��N~��,Zp Ͱ�K-b��n�S9Zȯ�-	��<���$4~|ΞY���V��8��l$�4���˸z�qV�R=��
D�#�w=��
����u�?�n둾�>��C}��j��3� ��ِo�1�C��Z��ʄZ"ۡ�o�%$��m��u��c����"71F��Ȁʹ�W�7���J���V�ī��ge�l�%�peRJ�I�� &OEU� 8�p��`I#����lm+�W�]K^A�K��N�6�+��,����r�h}�?��̓,!;����L�~��s�l�:�/o+����u����w��{/���E�@D��.�R�0�[B���a�w�4��Y\t��㫯Z|�O��(/)���H���h�좈�!�H6l�*������.x{�?��7�o��'��*t�M�?,���x?ƫ,�|�-_>�ĩ���_c�)�⑐ש����L���L���Ҿ℃��G�� �lus4�d��3[�_�����_�%$���3�Y���"`l}�,uŗF�бt쳖�ךM9c�^^4��~
7�E��D�u�_��O�?� e�o��ja�۽�y���@찊�+�B"���V�T���v�x�����Szea%w�0�4.[Ҭ,���
�C�K����ڏ>�F�3����5�lt��]�T��)��h$wiaa��|>?��D7�î��nR�� ))�8WO8���&1�n�R�vl������)�meo�T��|BPƔ���4����A��hṕu��˴��
�T��/��.�_^+��Ɂ@��q����ͳ��{�����W4�	#ހ�����5+TI��qqK]�h�D���'ť�-4%��m��/Ow�͗[ެǢ�6az��>�V~��a�Ж������Ŝ0*
�����ş��4���L�O:C'-8x�;2Guˉ�$�͟)}]w
��q����/k::�L����]�{��i���Y�.��=8��ß�l�珣��]�!]O�j�/:O�@�}��r޳uѦg{4��r����c���oj��m�_L[3^�����;���d�7#��^9*^�x���\M�Kn�Ƴ.��%&�4Mu�{�td�W:�	9�Tka9 |�=�O���\��I�P��%La�*[.�6�n�io�,���ɯ�����J�鎔P͌E�'�}�#��@���N͛��^�4~�z����n����z�^$�Tnx��P]����	�r{^�>���X��
|I�>7��n����d�#�۷�͂���K|����E�ݟE�5>nF�N�g�Oy��Ш��c�+�LLau��e��	���r�%>��Ӻ����?׷v���m���)�Q�*�Q�����Es~�lI�my����<~G�R��)�S:Xo��SNZ(�o�Fw�m�s��11�g��5mE��)_�Dd�|<<�ɢG:6X&`ݙC ���s��hi!=l��KN�Ivò�o,&�X*�.��+,�;�س�|hX����JArە�khaE��䗘�y�,թ�ƙ��+v�1E��L��-��4���6o9����c{.�זY��˳�o��B7yg�� l�4�O*SB���صQn���]�ɢ���rtG#ӓ�G}��R[� �²R�B�Ԓ�M�19�yyO7�A�w�RS$N<�4��NWW�����6+H�.G��@�q�֮��r��d%��Q=Y�����G�S�QU�2�����
IrY��FV�i��w�T9��8�2�Y[���
���m#mo���{�q	��2�6���T��4~���E)��B!f::aww ѲZϱ{ޝM�]���Ƽ^4as?�E}A��) dbB��_D���p����Z��HǾ�K�=��Op��T�]Ďէ<�NV3)���'��փWE��">��/
 h�E� �Z;����B��[^z�t��y2�=⵿<2���Yqm�!s)^7��w�}}� -u+݇0�b 2�G`jRZ�}�]�m�d��%������#+_�<�$Y��I!0JDU�v}������V�kv������W��h���h��/_�,x6�T���i�Վ�8F��w6_,m��&�t�o�2:^g���d��` e�bU�p�D���7&�0�<��L��ʪ�V��k+j��S��M�t&:�4z�]換;�%uN����&���>*&0�) T^9��͟�L�`Í�	`Z��߿����EW��lJJ����Y��d{���Xv���i�	����y�[�^��n[��+v�#��\`���
l\\\F����Zs4���%��Y��`l�í�<'�ud��bt[;V	dW�/ܢݞ,�ڝ8w�Y4ϊ_F��	16ӡ���G��f����Cw�Yl�K�[I?}�x��u6X"��%&&�	
�zh���N��2j�醢--\�a�˙%MLf�f��	�݂u_6��<��ߌ���uk4�o�;�oK�F���0���C=�=8! l1������`XW�����RLJ�S:*5@ۂ���H?۲��Er���T�!�q^�H����N��A3�F��k�<���\��\��B��T�TG�`c>|�-Sɳ�!�In���0
l; 柖�=<似������Qd������E���h��c��/��D�L_��8�x+���q���*}'�͙��]"P���v7ܐ�"t��#gr�|�pֻ�-}F`?�@_��Պ� ������ =K�35��#<`߁�OZ�����\_�1�\2w�.��l�6�~���d{#���08���lJ���C�Z+�l�,������=n�0�ox���0ă��a9�MXV
�4B��(r3ypw�{�����]Lq3���u���s����� �j8x�l�?��+��O�ZLNNJ䏬�~�Z��^�R<ܙq�)�/�����lhu�Y8�_t���ҝ����Ό�&ۦ�/�A�D(�����w�xV�#�1p����������}V��`�,�Y���[�����K�]nU��!���gu=�N<��v~-N;JotT�u�h6*&O�e�G��#^Nax����q|4�L�ݣ�V�����G\6��f��%�ϗ�([�x8�3�VH�g�6񪁮e~���]����m���:�N���G�b^��N���S��t����#�i2�R�B����P& �e+��~Ы""��\�2�b�_XbI���V����Ay,3J�H^1�l�ܭb�Ft���I!�s��y�Ֆ�K��)�9�k�/�1m;�lPA���"���6�����3�����^_�:���բ�����4��/|��7���H�_�ȝ��)�<PA�V v3Z�D�d1 *u*����HC�J�z�X>��`�K�RPb!���_t�Xu�PN��dƟ�XJ���仛�*!̬���N�=�}I�2����$�T����m�ભ�p�.h�$�t@{��4���\LU���p��x��UHDy�!k�	G'�;n�9m��g���F�>���	��X�v�.<7�`�O��3h����V���Mur�B�^��,��^SI�iɆ��Ɠ��n�M�*W%�>+ �/��-�ؾ�)��.dbB�P���1Y����j"�=���K�����8�	��	H�0m���~�=����G�^u���p�۪���Y$�/�IZ�\�D~��� �:��>Ƅ1��xi^CTT�^Q�#����vrZwiT�T�^Ky<o9�$��b���̩�H�VqZui��.yZTD���?BQ���RN7lβkc<KM����.+�z����'ՄQ����/�Ԑ��+���*,��!Px
:���H���INjk���q�u�O��L��<�t�m�����	����ڰ�N��Ӯ�tU#_8 �������o/����EWWW�CE^`��m�(�vޛzV��� �"�e���X��g��442��М���<��H�eҢ��"ٛ>���.((@��Rrr�g����}[IR��/Y#�1�l���
��O�F�T�X�Ǟ�JVtu�e+��7��S���G MՀZ�D���� ����.&�% �������nd�X��"����.�-B^���� ! Y��}��E ���*bb��X1J��aԊ���B9�N���g]\�ަN�/n�TTT�R����Lq�A���v\�}�F`��ݚK����P���!]� ��ߍC�}Y��C�	B�۞8�oC��i��h\�6�x<�ΏA��7�V��O�z�59;��wo㰣7q��w�U���9����T***$iii���j���ko��`�ɘ��ё�f"(6q�v�N�Iw���?�!��Ϫl�������K�6Rߝz��G8�꛶��w&�9χ�a�p*�o�Wxۂo���#��ٟ�g�`����Ⅳr&#��\z���0�0a��P�v?h.�b$���+>��>�-�lpu���*�5~˕�#V屾�����E��S;�!���@�N�A�/�_�r���m���ٝ/æ�3ߞ�E{�M�ԅ� vx�#�f���e���K��׹��e�Ow� ��8v%�����1�~���{�kf���̊)�3*����a�G�>sy��I=�*|6���m+�:]�fr�N�w�|���d�S�(@k�T+!�},K���+u���.[Q���jtǚ�\����Ũ�t=+�7`W3@�ߡ����k�s�F�G׏t�|-E����N�k�$��qೀמ��E��G;�:b�J����R�$����nC�۔ʬ��֊>c�>+�%j�p!X�����ƾ��;���}R̪z��u��n	r&Nx��ƕ�U�x�<`���8�"��������^N�]������o�3$%f�F��u�K��|h����G�K���.�����\^��=h�*pԬ0Dk}1}����g�!|q�ip�XY�Nm�u�l���@��q���P7.��]�'A�h+�s��>P��iX���w3330>?�̍�#�wP�m?K�`�h+��j��j�n��ed"N��^���u���OGGG�D^�J����Yۜ���VlL�;Eض��E��s��5�m/�y�D�QJ*R~�5��m���;��n���	S�ׯ3l�[./ף�Ձ_��?��B����u�(&���M�A7�?x��q����%;���v�S�8�Zq6�6��e�� 2[�4�:2��k���$ג*Dc�͝3m��F�������
h\Xs ��#Y[l��� �|��(D6M.?2��w�p"i��Ky1�`�7s΍�T�"���Ō�G+��ĺ:7C��=K�'4	fR��$���
W�ZGʃ_^
"P��4���{7��#��#���3�=W�sǆ�oq=�Ц��Y+s���qm��I"�q&��ܿ��bơbw�,!9{��e��F
�0�iΝ���ȯ������5��ll�"��6���bx�+O�"�sߏ�u��	�����X�Y���C�j(7�ѱj��C_�V*"���?u#�7���]�.t�$��L��qq��F��uZD��x�O���u_)��1�]�,^F
���c*��э�CyId�ݩ�AÚ��G}�N9O��"�x�L�KX�}e@�:�_��T�� m����8<�h�$�w~�
l��	��V��Q/��>9;�qz��9!�y~d���1G_g�+��IqͺUe�J�ԱCj��gaa���٤:%E�qQ���^)1qq�(���P�Sr��oM����e���A��.�N�k�8�N�y���;�ڇ�	=i��y��������U;rJ����������XJIC �DF�ݴ��?��il������;��rćZ�֦Mϧ�߭�=D�L=L&�@�HI��ur�gfS$,�
���e��g��g�FTWճ��<0�H �rVP�$��'p�@e�����a����K("�<�$�F���٥w����t�6.f���MM|����^�6�gS.�r�������ٴ\���c{~5�"r���
�������o�@6?]X��4FO#�����I���4��Zb��7��!Q��ُz�c���@muŏA���7�DJg�[�dɵk���ϺZo�l.=���ݚ������
v�K���k���X);/��p%[��f8v�:�W������:��x�����	�6]���/n��m9v��|�Y����l���J -�	l̑��4��F?�%r<�<d���Q�'�K<h�%3(u=���ͬ���Zҍ������p/g^��KP�k�����N:��o�20�����9t��t��C�g���`�)-��Y��v��h�_��[Qj��^�^�8?w��r��Jg��O	�n�Y�����YÊ�]fEfǶ������� VYq1O�'������K�g��Cw.�ӗE�%����g�a�gg<���� W�B�@HD���q�2�\e�m>��27 `{�A�q�3^������8�ʋ��F������'�YM��`Ӽ�1�5���E���Q��ƄG��HEM�p������t�kv��[�}�pz�μ~X��,LY_?:d򅄅�()�9�����j���':���/8�&�vi>���Zn!���?�L�]A���uF4Ow����l�h�[�vIZ�K�J��%h�Y�#@��a�����_=v�Xa&L<T��f�b�-�WN�����
	��e���PE $$t
�L��Q�A���ʍ���vd����4--B0a����	�v`���~���&�@En�k=�N�97���PȈ�䲻�[Jvdi#��K $ ��UUut��)���E��k�W><�X䡢�O�I�Q���˴adh�����$��Mc^,8b�_�<�^ڲ�"�kBw+)�����!��"M�>�0|l4Xm�j8[n�UC<�J!N^��J8d�8��Պ�� �����:��p�YJ�Yt�i��ڰ�S�	��xm��8{*q��ք���nB�Zx��jʎB|�)��xm��R��G��nGs�U�c��EDH��jV�� P��Y��ʷ|7�U~ϿG�Fo�z�]�e���4��m��[��ͧ{�=[q�������+�Q�"g�{^-�R�����=j��k
RAޞ���`�8��|k���O����]�~9����%�p�y����u��;�����Ґ��\�,t���t%�S�I�Rn
�/o���a]�7�/�JDn���]A�j��AU5([2:���N6�z3
}	ht�@,S��f��+�)^����Ƴ�vp8�Nþ�s3�\U���.p������I}�e��M�p��2���F�������5b>ʊ�L�)&de����;���"�M���~����z�� 3�;�ߒ�?j.O�D�b�*P���~�*p�1C��e�8�+����7Gs!g�.��#�O.,o�������]�%CW�qas�N��6o�
���`Cu�u=�\U�/�dK�5���Y�O�h0���D��a��j�u�ς8~N�!+R���UV4��h�;Ζ ��f�!�׷pģ/z���%��Z��;�u)�ɢ��ןQ8,3�L��{�l����AX�O2槾TO0m�Oo�b��W����Y�&��ك���������N��:�8,�ڑ�͆�VpOA���q�ǹ�[�T���6�`n�}�԰�
�� �IM]�m�����"��x���u�f����h&�']^��8B!���'�����Gf+��_�^B�!y#K�-;_��Ggj�����x��D��&Ѿi�_ȥ�l�_7��Cpxg��X��膵�H�������_�P��\�~F ���tH�y�%s�Ό1�TV���`�p���M�|H���v~zzzQ���<�w7= ��j�/)y�`�|�t"�����9��x�<��o����v�����=S���O����'�C�q�K���;�b�?N<��&�Ο�y��ͻ��_}�����!)%O'�џs�y��#��E7A&�ɚ�h�� O���m�B��T#}D����3��} ���|�P�On|o_XT*��4~"6�!	�'?���|�)�,L�;ЙWj�mN������
Ԏ�
#���t�Kl�S�h�F�{�,2���L���߉��-���`*`�F�ӫ��_S���v-�ҧ�e�D������]�m1]�ׯ �`bzz=�������Q�����mO�I��C��~g���?}�~��9��@0=�zzI X�K���]`��2� �2�tj#��R����Q��!M��x@��k����<{ݞ�!�pf-.1i���`/<@����{���z� ����Y�o�N�G)3������x�8M��)p#F�8�iI�p��<��5:�z��!)X�O�h�6��
{��
�3���#_��;�;.��Y��OHH�N��Sz�F�Ѥ���'��������cĢ�>^f���sU�������^�·���;��XCB�-��+�]������ʄ< �<����8�ҏ����(��swk^�M�0�|������2n�I1!������L\^�����s@�k�E����Q�r,�F>5�����/�ȡ]�adu�x��=W;��x/<d�H(�azB��GF[n�)ToP*��׵�K�h�Y��ECC#�����*�b����YP�RQ˴���gM��ka+4�=�\\8��"�E�+��8�ccX�z"�c�8	'��$rz��8M�a�KDcu^?w����s�&��a�g`����>�ʂX^qYY��i*�u�M�?�Q��]1�[6	fXs��8_�(}Rw>�]FC�<��-Ό��lh����� �`=I;�$�:���Ph���H�|j���yKrt33�����n$�6������6?�
�cC�n��|IQ�N�ujj1�!9���w!Q98��L#�xlY��ŶSl��G	�.��,���x��4��l/_~p�HPϲ]����'8R���1ɵ�u�4l7u;�E��u��e�#�VYj$iTEZ�b~X��]����J�x�&��T�&��WN���{��k��D�Ԧ覝wƐ@^"ة��f"�i�s�N�3��pH��Y����4��o/Q�c��/������,6��� *$��2�����$�RfP<�v[���7�Ӱ04��p��kW򠔴t�jg0B��r��{�?[PZ��4J��j�P=����2gY�=����=���I�K�B�)��0���F�y��FH�,46�����S�4�@Y>k��.�)m��i��_v�'A6>�V�a�t�hQXTD�gc	�#�p{�M@J��[[V(�pw胩�
����ދ��ۊ�(�ϟ?��,���ZF��p.��<��4j���+��$^��U���7�����R�A)���D��h�3�5�'p>���y���l�.V��_cد�d�X��/�:?o�+��qZ��7.��f�i-�A�V^Y�V�M�	�9b��$gd:�?R6vz}Q�U��ƨ��0�VM�S�),T�#�=�U�8���ٴ~p�s����bBU]7P��Qj_j�@�ͼW�τ`������E��5?�üR��,[�_+�q�%�>ҞCnq	H{h:?���3�J�oǅ��P�oLjE&��\,���G��F�݁�ݤ���|P�=����c�VUU�k%��ڶ��yݜ�������=�r�D�z-b�&�n��Qߓ����i�3���z�}�>�Z�
�(&!!+��"U L�2GwW�[��e0�%�;0 �n���~o��5�
��d� ��

z�m���X ����Lpc��q ��;J��8�ČM]��c c�;���	���|�l�I�W�7F��ݼo =:����z���o?���s�B�#+`��9 �m+��_ �k$_!��?)&H5��~4�ϐ:W�>��&KX���.����4�C�8�n7
�(�u����M�[L�ʣ�u�ط�7��<u~�x�g����,z{3����Ͳ��Φ�8�K>7�� �����pk�@��JS:Tp��=��/������Z��dqؑPH�>��<�J�F�]Ewjԝ8�[?7+!��U�������q_;���L�_�W��3�uV��K'���^������;��������7��ZuAvɹ>�ez���~k�(�/�f'��q4K��%���K�A���q�U��
�kh�})�6T��Z����Ұ-lm�]�@e32 HHHZ��ﾍ�֋��������&U���i�p�ݣ/"��;���h�,�Zb�Ϫ:?eoz	�t��=/_��sO�3#�$O����,��nl���`r>d�#k����==Z��=�D1x��,�J���n�:Ɂ��Y[_�p��++���RU�����yl��K�N��-��p� �NJ�7u,*��MZ䉃	؂���Q:�_�wƪ��>�������գ�չo�:v�H�=�.�֨89��������y�nP��g�^3!�dTW�����!X
��|�$22d�h7�l�$-*������A�g�Q�P�fo_7������8#c��6�����0@J�^P�<+J����2틒hs�o���ʎŜ��~�m8��Op�H=�Y[�~��~9*X�\����b������J-F:��s��$��}�<e��&�����|�
w���u����W��f+�k3~�Q@X8!q�]v��<�M���*����%�����S?uÑI� O�r�ɣ����<��ց�'r

�Ö������L�0�_�\�e��f)1?�9�m�%��Թ����d��San��N�
{�p*<��L�=��:@����yo�`,G�*���|�#x�U����
��._@��_��3u}���KO��g��g�y�>�q�H�hk���l-Sh�֑��]�1���a��g��'(&N�C�䏽o��d7m�g(x!�wˇYA��)M"��c�����2s��0��lG}���w���44��l_�,w����Sɪ��0�����)|���;��-~�>żˇv���	�)��;�\���YT4'}�x`r!�a�e����(M���p�#�[#�#�$9�
Y�_�U ����S�{GZP\,����߿�Ê��++��V��K�~I�2�y��1��:a�
�V?iV�`����?�=�>Z�Q��p����Q
��m�R�'�{Y�,���s��"��>��G*�iFW�M�3�5��wG�gڳ��h��43�(��:�t&$���cz��������Ѿ����z,�̯c
8����]�CI�M8H}M\ܸh#&!A�*�;�+����q�DS�kl������Z�pXV	�1��b��H~4Qb�дv�(!�j�z4"G�ɔ���ux���s��y���'A��9�Wu1۹�M��:a����������hE�Ta}���b�*J��t�s��ƀ5 �j���4=����
�*�ϨGQQ��?)�Y�ao��t��?�#�B�=�%�*�!(�y�qL��ڏ7ذ�w!׀x:�����2�P��+OzNo���A�|3�)o�Y��#���CL�f�m�߯����WJ��OQ�xd��Y�oe��ܻn(QΞ�7��B��Lss�,����H��3��M�����k��z�:����B�q��`���&��~P����F��G��>�])*i�����򿛲��(~3�]+�����L�}�e
<����5��Aڣ���OJ�UA0��E�!c�HG�2�5<�w�e���pwa4D<h���y��S�ߦ�oj0f�o齩�Au_K�Zo�	�m9��0��j��������k�+j�ݓH�@�q%cl|�G�_���9����uW�`�̛�O=�,��>�J���q
��sY��*�ip���(����ʢE�@K<;Љv~W<��e�n�~D;B����4b�H؃�\Z>~����R�����wu���t0r}�UV��Y���]\_(6V6����l����#]ğ�X-}oO�pd1�.F7}�tX���=v��:�}������x���p�����M:���e�a?PC���T��0-[g�M{3 |�_i,�����i�y{:��d*�8�Nd�ua���D����I�Z(Oa��QH�x��{��VyE5��C�M�3����:�/���߇���ڽZ[p²<H�4��T��ӲQ�1�U��̚�M��7z�N�B�vrCM�QT1�>-��Gnc���X�|�k�[A���1�� z��Fͻ�n�N؃o-�G���\k���~P����gm��贪m7���bюJ}�4��?��?���*��� �6��M�1���߆�_���be�S��� ,(܇Ue���Wl���mV�mA�+בڼC�'�<:~M�QS���7�ʨI�S���E%P�B
^�I�
��*��հV,���X%�iU!�8w�XT$p�is����'Ս�k$Zu��Y��kFo�Y�sT�OB�@-�����Z�_��^d���'��d��ɗ�w��O߇�����q2kkT�1�K�v9�uO���� ]<hF��m5G����cj4�n@RK>����Rӆ!��#�����-d'��_�覃L݉Qՠ�q�'I;�.oL��t����f�����~���n�@���Br�ڵw��͵������)0p�ͳŤ�p¤�����ZfL ��,(��
��;��hp����5�4�'>�������?��2�}o�O�.S���i�`��e��4�Cƶ�E��h�`���¾��Yg�W�Ω6&!kc�%�[j���1 �����Ńb��~&�����g	�.�_b�>~�c``�A�u�#���-��5�F ��9l�N���E�f�o���<3��Ϭ:;��j�{������~��fW5d�;��`�?Τ55E5�]:jjjJ�dZ-'?K�$L��&cy�g:���h�����L������� �9��E@p�Z\��ʱ]?�љX�x��ȱ��"�w�j�.��7����F^�9*�'�WΠ+'��gܫ'�g
��=��uUp�
,�:����sY]�:#}g���������Wu�OӒ:���N#��\�#\T,���,�'�Qa�[�JJJ��檫���}�[�����2��������N|Gw�:
"�h|�Rc'z�~���0+���c|�N�`�5�4]�?Y��ǖ�%�9�x�7��L���a�ѣ1��8l"���������1�Q���U��7J�{&C�C���U������[Zj�4����/�3�bbT&�_��g��s��*�|7��9���ۍy�3�;�1���r�>~���^Q�D���7bv��E�#��=B��G��{gvZ2<	$)i��";j�gL��P9�B�Jn�+1p�iy��?���'��j�Op�%ň���CB� 3U0ۆ��`rYl���W83����&I����S�[P&wd��z�����\n_-'L�/Ή�)�"o�u�
4��L�auqa�4�ڊ8�e��x#}k�I�~�s�"R(?i��O�Ң�b��m��LJl|4p��~�f<��hi����YSD��I����9������e�Q��X����C���-P'�7���<�S��%zu��"Wg?��Bw�ҷ�(���ɪbu�R��[ytb��7Xp��Ml����?� �J�i3(<u�Jǫ������v<��b������!��\�@7�L]y>0��u59��AL?����"3���:b��X� �~�^�U
��T�� �@�$�W���d��x�̢ڟ�H )���j�L��r���:G����ק���?N�v��K���l�<�]�i���oc�%!Vi�Z�����iO�
�}��"�`�~v�dwK�9\2�"��E�8��O�H����a5_;f�c/ Δ��U��.WLO��e�O��������B�����21^��q�it��^j��]�Ep�����Uq���-��6 <�z�='������_�>	��q�T�@$�@��9��^������b����k*��89���y�% �����_�@��K/�+��j+��f����2��m����aЂ����%	xq&�a��B���z����̓�ze�rrr4�����B�0,9�|3����LUVث����#T�����R�<F�ʪ*�\YYEp�����?E������������㧀GS̟\XXX���4�Ǆ�Q���۪�>���a���-�U������a�3�=���6���)�T�?��&�Â�q�k�Q���-xKE�"��4��
����vL���
�.r�HB.s�?�I���Yov]faG~�����+�J�\�ZXC��BB�w�� �_<.8����$�`s(��eMY��1u$ϊ�'>)F��͇+y�|�.�8 �S��"By����8!!� {W$
^16֮q�Ƚ�f3�?��A ��h�j�Y���v��½�*)��g��?k`���Q"�_U�I�(*�Mv�GBQ|���F�kT����,m�qʪ��$�;`�u}@��68�>��I� ��C
���#��~�܊�Ϗ��j�Z�A2����~��6�;���W�������=Új�paA��t�H� "M�tB��B�(�
RM:H/�C�P��;���Z9;<�{��?�:�+��Bv�̬Y��}Ϟ=CIF\~��963���o%��q�+d96>��*�~����%?%/�u>=��T4@򟅹�>���/�$������oQ��u�|�T����C�gwV�����T�Fv\IBހw�S��5�a�<a�!!A�򊕢񭙍�c�y���ӧ0j�,P�t�<P�$�W2� �Mhr�u�����z9%�����ݹy�������`\��bZ��N��D�	ۑ����_:ڨ��b?gX�vǸ���Y�K�����$s�{�iࣣ�t-�/@�2��.�A J��Iť.��G�z`�p�x"���D�44�w�N݋�dܦ!V�TP(��?�WT�\?�L����Sp>��e�Zqi���uz�޸�l����@r�2�_3��ZPk�Ov�E�HE����6Ӹ+�*������.*��cU	붎�`�<�N�����W�����n��Ħ���z{�{d��LbA�l�^�5�c6��~�.k)�O��C�)�E�^�0=j��β
{�<����H�W!j�`W��gV�\��S�Zab�ŭT��F��r��䗃(y��~T�a����"k����!���T�2=���({�Sc�|�$�|�
d��"�[C%��\k� Mx+����%H���`�����H}̀���yM��7��b��*��������"'�nsq��!��Wl7Q#�o���P"��B�����{�R��0w��w��Z���p��Ƙh�F���D�G��������]����׺����S��&~0|���b���O��U�~����0eߖ��Ϫ���1v�=~�x`��h|Y����l+A7�w��N��!��l@.�G�Ӌ�y3�Y|z/��6R�c�^��_b�>�_Kq,�U����x��_��Qu�r�	��������*�}2��-	�1	�^=��,��	��$�,kh(��` �"��B��ii��Y1���K����:���.�í���^m�8���������Zp��Y&ߥ���M_J^�Mc!�^MK�&�� ;�=��r�(����[9��c�f�}i�&M��E�y)}(��N:d���ZL����So3~�:�Op�G~Uf!�/+}���r��նz���m֔�K�q^}"���)2�-|KwP����UB��4� D'�ţ��$ �#MU�ɽ�w�~��N.�{W�%����ǌ�Z�h_oǺ�4�һ~.��T�ј�,nQ�~�po�ayC-Z���{0�Q��%�o╰қ\=�C���6�m�!~��]�m�%�����Z|�����9�]#V�z��$�b˷0�Y���yJ�T�q�wd+`����6t��m�G[QAFq�t}��eBh@rd���-ⵡ36:jwz��wPW�� ����lLU,zuE���(n
�9�K�����½�Q0b;k�3=3�b��r����n}K������FX��3`����W�g�o�[[��f�c��o\{$�Վgl2����{Mѱ�{�h�����0TnD�6�+��\#�?2��0D���hj��'�^
j5[�!g	Ȋ��n$B|Ĥ��9s5��nq��Sæ���/}]}�eC����M���^��^��Y���I���Օ�+-�3J�ͤ�x����Ub�͂�=H��Ӥ��&�E3���?� �m*��A��00"~���!k�q��;�;W�{�}��_�3	��Ɂ���?sJ8+T������iRST�~������f�9��j��������ֈ�S�5�?��/�8�˽|�����B}����΄<ys�Mڠe������CO��x��<��<�S[FAA.�$�����u,��_-v�j��Ϝ&(����x��0'w5$ߴ�S�`�薮ͱ�1egos���E^N�T;?&�P:R��>�%c�16G>1�\4K%�$�����=�����&d�Iȭ�/⁈�,��cr+��V��E��&EEEAs��FW� ����W��$�d�f<��A܌�6�+bHz#9�w�LO/�%��͑Y�P>����qܮ�h~@3��'�oU�w����h���
�Db6��{�|����l�����iOT����zQ?Y�G�L�~�U4�`ا��Fg�g����,�N��)+�5��c�X��"-K#��{N˝�sO7��k�����^���#>�̱���v�s>�VZ��W��Q�ۨ�Չ��xN=F
n�bmE����^��3�[�	=��gK�)`�"�ݽBuT�2.��«�H<v?<�M?��d�H!_��n2�Э�[=H�VJ�p/5���gE7b�v� !~�G��iJ\�5����ͭ��_��2���
�d��a5NS�F��?y�3�x�U�^Z[[7.AUutu�l^<l�bv$���&m��>��F� �����7{�ݠ�G��[�g��.�V8���cE��
�;��K8s"�rf���J�c�U��b2���S�١i���c_oh]�&�y0y�>=E����Eǉ���L�w�Jy8ե%ٸ�0��r�xܜI�ɲ�ZV��D�.9�O�]�#��B��kdi�vtpp!��FՇ�Y�ti�j{zVU~	�j�� �'�nŌD��%@���'v�:S���r~��C�� �Ձo��Ӎyd�-���J����q<jeY���e@Y��>��� j���iio_�Wj��I�ژ "�ǖ��eW��]��=�ׄI��w���ol�I�gy���0y��Q���S��+{z<���<E
�%�����9v�V�5_�ڎ�̸�m1�������]z`�ȴ6�������9����W"07/A�z����i/� ��N���;�o��S$5�U�\�_��U�`#���N#Uddd#ˑ�G���66���[j��t��Su��{8O����\�K�X/�'!g�u��|�ʕ�:l�a�g��wh�vƫ2��Q1|>�Nt�4�59��.��x��OY&]zU*s9���H�$�bڃ�G}+.��5��� �Z�"�ݟg�wF1x�ڮc[�����V~��d%UW�-����]���Ǫ����Q^w7,���;�\Ҕ��A���5灬�O�Y,�b⬻)s2�n��&=��.2ӤrU�"�	�9 ��8uq坦��~���jɂz���ث��C�(��r�6�it	��J�Z0� ;�W)����lh)��W�v���r��u~?t��c2�|�] �Z!�VUm?V�+����	��~�BqI�jcgɬu
'|���"���d�S驼�Iy�#�|�H��Ob)C
�η3���I����T՟���)��*�P�RA�i!TN�::7&�5��1�hɸ���>5�u����ɮ���N�n���.#Yn����gh���H�fƃ���;���|�%j vT"A���O���|w;h�Z�	:�X�S��똃��s''����Т�H�~�[� ��^V���I~�p?���7�L2o`b3��AH�~-k�cIw�1�<�@���v�� f#1)o�^���a��փ�(��xh��V�K�P`C�C����ɚ��E�K��Ϛ�v�J�˓�Q�Pݰ��B���%��Mt��Y��^�?���hjf!C6���8�r82��b����0���1��1""B�̬|o�=p��Tc�upߟ��W�!��� ���p8�b�b��iO?UQ����х(@���kYh���̖lU���~`�&���]��ƈ��ߢB�e�Z^>K۹��a�Yot ��OE���?&޳^��s�b4�7�4M�c�R~��H����!��|;O�~-u���N���ap>���M��pL���������A��{���%�߮��U1�1Ť;�fql�\�d���n��~�ۙ�E�i5��ȉR�O��È��F1K���O���P8#`OY�p��G�QS}�56.�,o5�o��"5#�� �]6��Mqg�f�5wC�����������ݗ�Ci���9��c����h���嶠�0�d X/�Y� }�xٕO��j \�D 4��9#��陳���/_(��6�R�Z���d)��_Y��V�����Z_�vީֹ��(��qE���P���%^�����,#�b��'�a,bC�<�)��q�'��g�⸭jl�^��KZ��J�{���W����#�%�U���C��pe'�Q���t�u�58x�U~��n��w:�q�t%�\��<�c�l��� ��?��G��s�l{Ӧ�^�RlF���Bj���ET��P�9�j9o��0�!<���IKMMM�Z�n�3���v��&Md�gA����A�[JA�MR�_����z*���1���r��}�P�sd՗ڢR�I����*�}l�
�$�� lCgھ"+s0(/���\
0j�q���[L�m����adܿ�����[y퐨��/���lq��N���\ʂ�6ZZ�SR�n�r�@*1�w[<8�,�Z����d�V�N����k���� 5�7h��PwrKV�)9��1��o���(��j��3��o�M�0�St�>_>��(*,T����䫧;l�99[H��{AMM�|���7���wπ�Y@�Nh!;u�N֬AGQ��KY�F�+9pHD��ણU�Q��[U��e�-8��Z16F���f}���>C��M���pJ6尰��"��ï U��&l��Q�\J���q�RH�h��X+��(���:0�̑�G�qh��\Z�{�Q� �7�^\����@dg�A㓓���S���7���
�~�ޔt�K�b�U���i��C�%�OAzTk3�����x�s��R�]��.7m�\M�� <��5�SN�S�?JJJ����a���2�� k�@,���p3MI�N��[sN[�g(�Jޯ��4q�e�
�����4=Y�d�P�U�h���j���׀H$�Q�æ��bS�#�_'C ۈi���8�r[��r#�:G�������@Ds�E{8'#�G�����?9��굱گU����]���b?�D�\�4�oh�G�S����ZM�\"\\F�WZ�Z���H]U5�Obf$j�9E����]�~���'��
���֖��7�H^-6������NU���אs@O.�yi,�Z9���_�n��j�O��Z^���Z�A�n�y���_tl�����U��>��*\.�u��^��Xym�����NPG���M֮������dvK�|L��^0F8���v� �dIsX0�Bڭ����t*���0C�X�B�j��{����,+��=��n09!}�[v��i:/sܜaRY.3�O�r{��D����-�DzU\R��0+O%�r�@C@���SzI&�j��p7����i����k�'�=$��-��a�Y��Nw�Q��?H��|��E%1�W�4Ⱦ��
N�5��Й�ۄᚤ��n�t~C�ˀIbj'��ϱ"�W��9��m���h��(Lm6RU(��+!D
r��"��~�#}�S|0��c���ax� �fS���
I ����ݨuF=��!����ט��VE�h��7)	5��d��i�F��$� C�,$UPPPض��/S&8u���.�L!�\e5C����}�Ky�/ݭ��$�!݋�K�hb��E��I���k`�&���3B.sG��V�����t6KMG�ƨ�*���c�:�l׼[q鯢�"��hM<�D"�_��wZG�>�q*��^�;Ϙ��f�o���4���Y�V�p������L��䫉<F�����	�ƽ�bNN��z*�unO(��n������etR��7�2���/��e�#$^���^u��ߡ�� {Q�P#.����,�@POo������؍����u�(hq�Ҿ��O�Ρ12���#|���ũ%������gM����<Eŵ�B��!u��i#��4�vZ��F���k왯��i7��g��ŵ�|F�%����H/ r4�m��o�R�檒lR��dY���2�����B`0����

a���b�!Z�D�Kl�8@xl's����?b�&�'Mv-Ҭ?SЪJ?��99^T���'��'Sj�(@5JEuO�wY��ɠɈ��zM��;||�8���<���,�~�uX���F�z@����$ww�˱�!�����JHH��?j�Mq�{��ذ`嘕d��eG �	�
޾����r9����%���7[=�߻��+x�M	�/��:��g�2��̾����?K��v\�'P����`���cXgP���6qʘHצ���գ�L�3�0
?��TB�gV���ڗZ��xwR<��?�����&���.i>O�h1@�0]���{N�;�(���X�l"���a.�4�ݓ4���ӿ^���Vt���G�u�S@ �@�J�H�'�����I�����4>T_E����׵��c�/�zs.���w�g�~����n�C.3a'\G����;]#a���~�[�m*� ��/��O�g����G����
9�KZ�\F�\%�^<k?�m��Ztpp ���ق���wf)�I�����'�(H"�L.+�DI��7�<�b�3���s�S!�v�<e?��1^���;���]��){��rcGԔ�,A�SD�8k����BT"�ӹ�e�OWC���_.�[�X+�Ŗ��/��&��%�Ҋ�T	G�q �;�c2]D(��틋��B۝�X��~l<ۋg����I�{K�Φ絢I��蜥#��=44���	4�A��I[wdd���W�cm�%�,z��KbR�ګy��dy1'�h�>O���s���{���/ٖ���t\�Z�N���������T�u�  f�^�sb���L��9r\go_�>���������Ykstl�St�\�0�'� ]}8��H��B�<{j�ڃ��7��j>�=\?_��t�g�PƳa��k-^)v,�5l<R�٥�$���A_#T�{E���� � jal�L�-�D_Na$��fԠʁ�S^K�]��G9|��aI~��8�myy�8��n��Bk��4F�(����B���7�����0�"��G�S�J�I���-������7��)?Gka��H���88�v����f@q2���4Ŝг�ܖPz�^�_�L-m�{_yx8O5�T�e�/��c����uɳ���R���%[��~���"�v	~�7`'�m�7h�t�����9��%ԣ��@-0��������ٜ~`3��ɮ=ߡ�x�!S���Ed�X�j���4��7�8�=��O�|^k��W��%�|u��8	�ee����P;5$&�n2�q�%���0z�oM�mM}��Ժ�T���3�{�<�O�Ƕ�B����s�~�� h2��wмX޷y M��{' �*pri�&�T�*/k���:x���J]C]�e�!V̶�Ntv���6��<8��A5���g�#�\�e�.-� �ޓN�n�f���O�M��;M���W��� ��&Z�%,�b/}��phej1�w�������H��}A�`>���m���7$p�%�Ml�m�䷖#o�Ͽ���T=%G�=۞�
C��Q�I=�79����-�����"���?n`'�&��B�)}��AAKK�9i3Vc?2Z��3�~E|�?.Hkj{�q��V�'�m�'oa�1�Ω�*3���-��
E{��jz��@j�YF�|�q�J~��'6:��(��� �Î���$�S��sj{�S�>����r4�j 0�z�y�5"2���C�j�����Dg�����Sy�F�p�aZ�p�":N�Pȃ�����V-~�kJg`��"�n'��5��]8�>�6����:Bw��q������t���	@}0x��On�2�^I�u1���[N&BH.<�U���g3��K�Dk�$��F��̂�x(��Ɇ�R��ۂ��\'_s���$����0�H���wv&oB�����ly]�xf��y�J�q�l,EđqV}���r��kk���g�HՎ�5�/�s�%�83.��a�����W��]�U������Y��?W��ҋ�r��n�����M�::Z��`5�5Tkح��TL����I�ۊ9n��Ө�󼜻�Yx+++� �\~[�-%�E�І)��nSќԍ�e���jk��<�|�f�����ƛi��T̹��b�bY墢n_T��I��lǴH=o�������
�i;;;W٤����-��G����$�3�C��yW���w��QG��-THT�����Ŗ�Z��z��ZUi���Qn�E���p$
p�4ٝ3
yz኏�1��U-���j�Eo��A������$"����ҙ�-����~��2E�0�;����u/[�)uM�U/&�lE�=�8���e�����ΥƚkR--��B�J�speߞ_&�I���/�&2[����U�^���$�\+}���7
������9Z3�<$]}mm���5+�9Rg�Į���գk���B�L��c�[���U��
�[.�>#��%������k�S����}uu�ls��X��!_��]_~Uz���pF��z��x|� V:��]=7T9S>����%�<�'C�bf�ҏ���..�\"a���MsoO1�F��.f��R獅E�-﹎���@X?�)�`'LaЅ��x�UZܭ�0�9��g.���K.�r�����u���Y��x��a�ӫ���)2?}�G����c'��
2��\�(�h��m���Dㇶ6R)ܨ�8��e�5�.?n����m�&^�z����%k����Q���C��Y"��
;�ݚ�yR�c�B �����(����.�4/9�o�{�9�?���)�ۦ�\��8e#�W{�f�$v�W<sk�
�,�-��98���R0����T|��&;@:�|�@!��,���~��U8���ڇp�F֋�H����;yI2$��A�ߺ������C�������EY?���hq���:���4�!~��"�b����;+���>'77�]4�JG_U	6=Rܸ�W\�m��(����p��c@j�+(�z=��{�:(k��?2d�fȑ�<f*7gᄁ����-����}�o�E�kJ��NN�N���8�V�[(: �MDD�]���u�&�Nuؗ/_>�w�}���볉��ٚ���
9or��M88g��%�j?��tl����[�]�����`���
��L���́��R��,pG�_���l#�*��4�M �GgF�Gv�CAs�∗�I6��ܢ�,!��m�����=	 `CqQ�[���KY��;׮���f�j>�?`9�������A~�{�\�l��M�Ű}�%$J�~xx�:'?�Dx0�3�e�@� d��8����?`Ap�K�s�Tb���LК���M�Y��\��;l�X�2^Vm�\ݷ?(����9�СZ�6�UK�.��sx��~�Fm��6�~�(:)C�dP�]%w��DG�D��nS �QkRb��b:��1�Š�&�xx ����/���f�B�邴��(76���J�z�R��K���wT�#;������c���Z���*$&������(�9����T"0Er땎&��.zH��?��/!H��X6<����aiy�a��Pī���pT����Ç:gT���T��WQ*;��.�f]���Fupp�zZ@[w���P��f*�����Ө}���k轘.����G�s	�faad~��%l��8�6��7	�����S�7�\�������� ��2Ryb:x0��0'�a6��12*�.k|U޺��E/f|4X��ç\\Z:|�Z>��i��s0�O���MBs�R��W�+P�Vm_�=���"'&6�-�Ѫý��|i-1� � P@	*mVg�j&0����Tjf�Vtv�|G��'���'���8�̫c�v��h�[��8��=�0§v�nq��m�K|��햟�9�l�Z�Lp����k_CqdTl�dd8������z@�x��$@P�΅,�Սs�U;Y��rQL��v����Al��A��dv�G�]d�/~{���8j�Җ�JC�O{y�!�oR>�yi��x�*�$-x���P���?e��DKa$�'�lG d�ʂj�#|-�@�{��8ߣ%���t�ZR>X���쾋�����jp�	�x�bV�Ƒ}}C��f��]>�cu�a�x+%���J����!��d�MГ��/ͪ�z�xE��_�
g'�R�Ŭ�8J�,[8�-��ly���r`� �������-v�L��k��N�L�O����R��	��{�FZ���Ơ꧇V�� :aG2�|b\��m��R��ls*O���z`�N�lZ�4a������މ��6u�}���NS=�z�$ڠ�x�[�r���+0j�_:�]>�`�lm�?̑NJ��ic��r7���u���"�WW�s��剔�Y��k�P<�B�r��|���~���uW��ӏ��	�8���ƕP_��&���O�0��=���ɩ�����Ĭ�j�bD5q�C?�7__Qh�a|�6F�B�P4��'$�!�E���	��{}��q�"���]�r����j\����G�wZ�UqƎ��n2R�c�χ�ʧ�Q �@>�C�$M����0��
��f�kW��>�:$ܣu��ע�.A��bF���O��s�(���l��m��&q�i�GY# N�D~��+���yT�`P�MEE|����혭��\�kd:�l��7���{�pl� �	^G�./�A,���n�(>u�L��} �� �Ԋ�Tq�rm��VG��\v��{�Z/(^4D�|�������pǈ%�;:318ڪ�c�˞e��r�s|Pk��2�nI���fl�.�ztG������K����፭>a5:�������/ZxH���Yn�.ٚ�&�a�8�~)�r��f�j͒�  #(6�kvZ#@�:�]_��ه/KTD�(`�&���t������������%����1����/5��)ϻ~�ݖ�ho�R��17L|�3�\3uv����v�6a
\��ܜ[�̠X��0m^b���w�Za}��ˏ]����R�'E1N�U�|�3	񼒠hsf3�4��9G�N2��IOeV�.S�+��I'���a .��p��* ��䂤I�� ��m�IGG�/����Ç��hb��L��C�c���e,�*�����:u4���s����9�|����$/pS99,�����MwLHVV���(�h�`E�� ��YP������N`{�Hnmk[RX1G����;OK�����o￪�4d'�.^i�Z:�ܐWB�ڤ���H���V��ӫ�$'� ['F����?K�#;G� e��0I0���7��U���=go,���vk��sgL��+}$�������ɬ:L�m��E'3�����AP{��a�s(�wKp�%W:�W	�x���"�·*���U��c��I����m��ۻ�߽s�V3L���f��$3��ʯ�����)��c��VMۦ����Y\H�_�9uZ!ă9#�O��yl�ds����_(x��7 '���F��>R&�O�P�[׶��f�ш�Z�Zm�� �kW �/_�~}��{kܟ��ă��
�l�"bX��2�F�[s ,2����E�1�m��M�΅9\ш�:/���G�i_�6�YTT�з]�)���dg5}q����:�lqo��奕�Y�$[��넻��=O���G]��REwn�S=�s���(D�AVoo�	���c���cZ	�T �oF�V�w��Z����ʜeYZ	�֊�G�Ɍ�]a���/?�*�����i����>*�<*F�H�NNf��K%ʞ�U�ʷ����e��쬠g`@`�STt�+6<�jX{_��*���W�/.G�mE�ZFt��~��RNy�rOO��AIYY���m�	�o #��Ck���&�FF[Y��u���XY���?�:88������ɐ������������g��&fk����X��" ���;��xh�����j�=<�=xV���"����(��'��Y>��f�|�F�vl���8����'J�J+5��_V�C�.5P�a=��Q.%))� ��9ݑ<-,,��� s���5F��c�8Q�U���<��<���3:���[E�3d/��z�{� ��z�^v�ú����pU�wQT���H����LD"mZ�rĵ4q�V\/��c�[�����o������؁\���A"��p9�1�a��@�?���6�R���f��ȧH��a���_7�c����Ĵ��:�q�E�WtTH�A'�����"fC������Ծ~�ABѫ�6z�gҙ(�E%��`�DGj����kǓ�8hi�B�괃���6�F�:Qa� �������lw���x �}d���|�96�ў���E�x���s�bqy9��9)����W��
u贈��S�~�6,���!�w>�����!K��"'}G��?	�S?b%J������2d���{�J�$��Z�b�09�i�b��c(��s0��M\�����`�D|k���������7l����$�渋+�L�>��+�l�5Ы1�3iQ-($f���z��R��p@��-��M\��ޕ��-��'���n�n�O���q/��!�hC�*+��2ɉ��s}$�2
�~/cL�c�|AA��e������ ��Ը_�X�`�������g��$R;(��;sƭ�"������!5K�Bk<\":�N��Vtk�b}���}���3�ߑ���־���d ,Y^Z�편�V#��9��/B���ڧ �占>S�j��o\%��@�x��$e���"V�o)���v�lF�ι�&&��)�h��63a;\�rb��x�u��a�NDR�SP���vCPn����U�P߻G|'���)�|�z����.}� ���X�
�K���K��ԡ�����/,��ה��u�P�0�Tr�&&$�=�Hw�v.�u���)~2ז�?�p��Ѐ�����2AM�R��uվ�6RgۣG��9��*�]1޹�U�ȃ��l���B�Ќ	����=��o���-���`��DkCz)��{.�]z�����IģJ����G4dƪ�7eE%H�Ο��y2�)\�=�B
s���lyi���u�y�ʦ���?K����_�]��Mv!�Z/�e�l�X�K�~c*�P��tK ��K������.�*֐��b�I:�|O�0�r�o8����BИ�iV������`F� ���8�,:�%k˴�J�@�U�P�zo�|�8�a����S�"�:"���c�������$3>d�x�����F�����G �OJR�W���%!�[[N�#�Սc��ƫm��]<&w���5n�� �c���ָ0��W~�cd/*,|�K�go_t�.ٳs��S�m@�8q-��9^'�e���`��Ogg3� G�B�}n����_h'�=ˠ���,���uw��;=uM����nN�$�:����#���Fbh�.z�j���#�xz�U�(�@Yv��o �/�^o<���.ś�s�z�0��brgխ��Z=�:!���K�'��?)'ރ�B瓬O����=:������=qR���u2��גv^�+��b�[x���\�
o�5gn}Bη*�Unj�GS܍�G8	��e�0[w��I��I���W�����m{t'5�{���U��`o`�`�U�<��Mެjp�|�x}��UO�𡬐q�5ܫ�� T'��F�]�[�i��MIr"�97P��<��8�ՅZ)T�,s^�П|��E�Y�:iN�x���J;D��1N�t*��T׎�:���LL�����&��83߬B�x�<S������J]�>F�}�yU� ug�5�bM�#YT��S��:��>��P��V���z7E:ß�1�S�J��=��\�W;�p �ז��}�{t�`8�=S���h	�i�k@!�[��І��v�=d#�!��셥�,>�h�4f�vG�}�E-ܪ�c27��]Hj�[�5������d""�0�=�,^[n�;O�9���N3q��:%��-F�=���~W��� ��3��/�����f�^�^��43CA�Xb<�<�u1y~�RR���Ma�n�u�<.�$�m���������V%����dzԢ`�e�L9`8�$�:a{����RS����WQU�G���e2'-�?�2`Uh�;���+$ɄfP�H1�j���p��C������
[� ��Y���G��ϒ������+픰���/���R}lO��9=<\0[E�wkL��g14�
?&�%G� ���8GZUՙ'�/�b�	O�%�'�Q3��j����'�/�H���R2`�5�g��:�Z�JoU�F-��q��ԓn��[�\�� Qpѵ�H�\���ziY�)�ɞ��pn��a�٫0��c	�CU흴w.�m�� 6P^V����n���^�S�:�������!��KxF�:�������<��k��fV�ҵČ�RYy�Ό�O�#߅tD$���
y.,-b1�]�<yQ}�oL�0��)rN�Rj1��������YL�[�� ���l�����\f�]J��lͶ�G_?}�3�^�?��ݖ�����E{PI��q��쏯�w��A�2D�YUZG �y5t�$��*$��c؋��6��k���˴�O���j?/�oY9� &F3�6�;,��c��M'��M��=!�r'����鲐J�D��������ۃ#lY����i�";�ϒ���,�C|+���|xZ�[�9�|�Xw���tl���᷵ۅ2�Z�_���R�6��4崞-�;�% �0y�,�o����Zy�!(��5��o��v�|�������e�o�"��12��4��3+ ��/CS��	��wfAS�l�S����ڎ��q��z7�TG5��+L�3n��qc�AyӍ��&������L���˚�BvY�J����ff囶�NLʍK�"�~ؔ'%%m��ϟ����\��·�c%^GRGl���f���a����z��Ve״q����x��n?bg�a5��6޹�X�Z�oX�W����im�k������b3̣_Zb��h�;S����}A: �U��?iY�F���6Euuu}�-G�;�/nX����=*�L�ՁA�7i��ѐ(��${<���7xr�P�=Ç��ط��Ɲ�S|֢�7�%�頿���'gv��oH���EC�A����9�F�T�x�PΞ�@H���.�o��v����t�&�02�M\t��G&2%?�o�Kb��ߧ��H��}�-�@����0��PB�m7�r���6e�9�ZeT�\��q UTH�8㲊���nmbϻ���٦K<1w���+k��1&AH�,��(�����E�kZ�*��Y�V���E��U_Ma��]o���8���H��
���&�f�ۄ��	�#ο�i��Eˀo.H����e��s���� /*�3��{��2(:��G6������ �HQ5�ϺmG��,����m�����*͕���������i��ߘ���
��&������˄�r(�=�����,�4��a�@F]N������?����I�,�bH˯)iNbA�p�X]�I�{����:�a+�V�
���q�<��~�,qݢ��m^H��C.�EK�X�'<Rc����߯9�ˆa@�ͮ��?(fz�T���6"b￳{��,]3r�2_["D��eee%55--��.�1�����#GF V�?7q�����&�u���d5W��1����E�4�����;���
�Uu��f���](�xH�+"5�6���g�c@�֕�~�ꪪ���W.��x������x��5�e���D����L�+օ��1*�G���/T.C���6h�^�������v��R�^��×/UT"�^�Rk@?��NЁd�f.����݃_�^�����5���*�D��*��dwp�=�S��z���C9̭��G@<0�Rȵ+���5mb��p�̬�>��:��^�Z����߁]O&��hV5�Eo��ޛ|09F�-7b�QT_YY�����>�g~ҹ�����[U��a���P6��O���pO�}��ļ������o�6��.Zf���D/v�aK�v�Z��T��)+ԍ�)��Y=t6�vӊn3mh��<޵������U�I�/����3�K���G"� �b&R���jG�v�������l_�T�n �Q��a6�?M쮞���q��1�A�Z���A����λ{��r�:>�So��-+���ƐD�<L�`��gs���gaa1)���g:�;����w�%��W���~�ġGo�W[**�1o�SN[�#�o�L)\�6=���s<K���յH�^;��⺎3���*�)��wDx�C�؝���Cw=s�
�!~|�E��h��d��U��r� 1tl=��l�'�����8{����0�����l�0���̌��455U����OVYG��qh,f�[$蚚n53>w�DF6��wz`v�? ��ޚ|Q�#�-3 �-t��]c>}k|�m��r��˂K���9=gm���J����w=�B�Y/B���r9�)����o38�?�I�d����5Y#-���!���n��Ԑ�ij=1(�Eh�Q�@\r�ݢ:s��t&���:��Ӂ����|����9 �n[�O3����G�)JJ����̉:>55��M�/���ё���q��?�L�h��)��F�9���ܳjx�u%>)q��w�%�F����Ơ�|�ɢ7���8���2⡹Oq��pڑV��a]EE�uo�37?��\�ϯ�w��c�����y �Ŧ@��v�Q����-�����n�@O�ҡ��z� ;�&�'$���Ϸ���:SL-LO�w�i'�A�a���%r*��n�;�]���w��Rd	�:R�19Ġ��_S@��?��]Tg������J[DG�C;H��0#�ۓ`CE��- ~�=~���2���:�3� &j;���p{*Tz��������[uٵ}�(!����4HK�4�t����t� �-H�4��t7HIwK�;�u^���~���3�g��0�#g�s������u�
��E�J�<\W��,ǝ���P�ZO��%�4)�Ng�7�*ʆ�_�45���'k|A����q@�PP��$OOO��}wL~��r�}||�rGo���k�3��FMp[V��A�}A�v�+�T6c���j��W>��<�P����Ef>�Օ��̫W�ެV�����;�s��X8�0ɯ%��+i��TN�����%�}����ȗ<rG2��~ٱ*�ƍ7�K���mز'�#/{o�S�*�������/�\�"f�F����r�n6�3K]��S
R��ǿ8x���ʗ�"���(.f���~& p�PJ�ܭĨ���w�ݗb�8�F]>e�F+���N���&qB�--�����e߭Q�1�/C�|҇�O(ͳ�em�e�@�J����f(8	���9�@����o�I��|�_�[���a��1N���f� ��OU �ӛ��W�(Z0�%�Q���Zg%�����{�ω��_R�i2?x�0�Zc�-���s��D4�h��Z�'1���/�C��o�Ds�ߴ��`�%��vkD�!�	mQ���3�y��c����`���ٕ^ǞS���uU�O��d*�P�a=��o|�%���U���<�6��t�V�Dn��~�˥2BV����:���u����?�R{��I� �|;��@&b�o�z#���sfɽ���	F|��*�$����������3ڳ�\먱�y��sss�~e*L�9��m�3�����.��/�9�ڌ�Ri�m��� ~�bL|�W9�~��*k;���.�mZ�섌���?�gN�w�m���L�R,l��Ψn��o��9 k�k�?��v���21���tK]
�+)e^5&���9+�0��<�6�A�fX_[�(a��g�����"�@�D�;��Mi֫�f�볩׊WJ��@�{��c������d�I�Q��cG�	�ؑ��'�G�5�9r��a��T̼}���,���YK�=srQ��;���ٽ.�/c@�`��#䍢4�9�����~�.m�RV^��{�Clݠt�p��{1=�:J)����x ������2֣���Jϟ?[�~�~kR�t��k�ׯ�Q�n��
T�pO����f�����dS֔���x����y`选��ip�V5�D/j����c.L�M%zZZڜw�ZLHp������ X
�5S�댴2S�:�	�]�* jo�>�.*���=�����J:�d�v�zxtt�v�j�0A�b�����y^"�ʱ�P�D�_����Y�6��~~��B������Fg�;��R7��x�W�[�y�}�CED�*��4��D���x/˚Β�%^�����3�:Tɰ��T��!}PG�{�L(�ĄI��C���cp5;s�#u��o����cފi��Y�w׫"Q(�@���Ai�6u^=i���s�Dj�zg�� �x���?���p����pn"b��@�s���`K����` �*�*��7!���t���d�52G�����n��#����q�,�hj�候�����3��Ic@a�Ȥ>�0Ʊ���Xl	�\��1��g�(�6u�E�Rl%>[^����+6���	=���˅�(��8c�lɩ�V��?1��v�=�U�<�l_�p��v� h�s�T������+K�f�Jmj����?�����c5Բh�c�{l�\<�l^����J�ߔ`7�;"��ˣbdD�8S�i�ܿ��-��K&E��$>����Ѿ�]WG����/-�z�����HII���'����!�2�N&�8�S2�4*%��ۤ\�1�#���l��O$������z9���^���-�NWL5{7/�A�xy\m�������|#�QV�9������j�yIlju�
���.��0��Ey%'g����c�p�ԭG0��]� E��^K��8d?
2$c����-�a����K���l����f���ﯪG15^s펯�Hoߢ�V���S黻�f7�B���2G��׫WbFF�F�Ơ<;瞈��J**������V����{ �n8`���-,2�+?�5q�w����uu���*X�����������!��?�-
(:�6�J���b4,c�V��F�a���l~KEkp/�K�4ƻ>�&��FW!�;F]��0��3������;�G�R�%
X%�hz������8��vu�b�$~
��q&������C@�H}�� j���HN����63ζw/Z�Z��Dc��,�/�}�����V���[A��N!�%L�,1vyjJ���#��7�� w�@Ʃ��i˞�~q}}�c�!���X�^k˪`Wj5����BΥUߌO
�>��>�ox%��]̗1��H��jR����o�tY �F���|�A��A?���t�@ȱ$ʕ��rE<������!	��2��y<bE��ԉ�ul��d�Sd6�nN�3Ф�GZ[�RpH�YU_ߘ��ڄZ��m66{��'{�nu��H*$%hSé��Wݽ�ˋ��'_���$��(#P��Ж���Ԡt@��F`��	A�?�7�h5�( 0�Y^��9����TO
~���W6X��?�6�l>�=\D��-b�Eiu����{v9_���4�@[Qt��jq��T<. ���z��=��l��B�a�/���VQ��k�L�Y�����Kƿ@�g���%z�-燬88i����(�>T���UA����@��/ٸ����qr�<�_X�2rv�3�v"|B��-�u+F�L����W����c�*[T��DP��~�]@*�m��
�6{�|��JU .������+�0���@j~��p�+�j!��z:�9 J�J�?�?!�v����r������o��;�Rx�	p*��^�3��'y���d|��W�'Sg�R?}k��۟��D_8R@
�/��|�wo��iϙGi)pz�GC�=��NM8�)�f��qX0�W)��dr�<�t�\y)�ܯ0��/�+u2'�>��G��p�%#6Q�[�q���J_6$p��.�D�����%��{�*Ы
�ES3��(����m������Nu|��h�������
Ry�/���#o���%���Y��;�"(�z���``�z�ߞ:�����Q�2��籹̰mHؓᇑ����T^I���Ư�����\8���?��pd�fL����#,�p��Pw�1T�����w�*Ķ���1��ԘBr{YƇ�h�P;��g��|s�.����O�q�O_�o�$󢰃~����M;�	�klz_)�ЛY��bq1�^M���,���=��O�oн�]�Q�����E�߸U�#��|���OMJMH�ʤ���~ *ǅ%���_�5�&\�A����Q�L��!�A{��� &>�z��+���٣�N�O��]S�gK_��6�����[���0�x�����.]����z�.Vcy��V�g���P�{��G����$�����'p@��m� zԿ�R�<�[�,8\���K3T�(��--�*��ä���ږmZ������8��B�]��H0�$��<@�{���)����NB�s��б\�p�;�>��y�絒t�%F
����I�RO�������	�����Q�V�,y�Y��F�ډ����%�ш�!��a�R�O��`.�I����Y4��!AMC�jT��������(xo��hj�
 ���R���W��
���QUWϪ�|BCCCn`�k������hĀQy�%w�g_�+[J�-�F�s���⒒���	>~PE9L�h3������5A%������qN\�/ZU�[U��N�9���e64�b9�����0�ʉ�D[����a8J{W�a����/����[a�۾�/}G�|6�zd���|F�0J�bTZ͗�*!�t���|�"2��ќ��n*�q�ehcQ������͟��sebf�����Yɸ����(�i�t�m!Y$Ꚓ �e#\�6kE(�K]@n\�{�����~=e���gu�oTT��i�E�qζ�>�GQ;�lD�ڇR�pa֤ ъ���ۿ�yv/@ǡuω1��%���T��Tѧgf#����8g�㵉J��S���|[r� ��:d�,[���{Q�Ì�[:�O[�rD����B��7׋�R���C���'nB����ռ<���A�����tk��Ag�Aft�X�����l78�T��������ψ��<rמ�*�
�e������e$�x��Oe{�2Ƿo��<pk<�`t�������s����Ov�V�K���D�Ni=���N{3�k%�"##��.~�Vn�=����X<���,�������f�vznT��£!fM�����t�!N#%�g��z�G������W5b���Բ����e�;�٣�� �|ym�dgg7��5�A�(H�V����)Z-޵Ȅ:��6K/k�+�9�rrs�����)땬D�IW���î�$��"���o<�v�xx�VC�aw�����/� �I�S��@���r�OI&�2��������� e���)�`ls�'�hм���Km�����~(�IEm4���x���.G�-

����'j���Ecc��8�zᜰo�է��0io��MR10� �'�dѫ3l����a�*Qdt�lȖ��{�#�j�5�,j�2j�DЩ`�@(rD����&/ �w�˘ܹ�(T+��u7ޚ,K_�U/�y�q�����w��s�((	RR,,�0/�=kkkR]

�����,�C¹
H�b�D���8T��N	�RB�|��}�����h�/�۴b��7G��t���P���mk���C>mںJ*���0*�-���f�j���C��M]���,%Ƴ�S7����
y*�=�� 甔���~���]G-Hfk�U����y���V�f�ک��Ty6��Ue!;(V��m#�������^�������P1�+ @:��O��g�(�x�  �w��VL�'&�[�H���1l.4
 ��S\m��W�.4MsE��să�N���>ø��Y��0Jc��$JF���r;i���}��B-�`��\ ��	��s�=��)C�����;����itw�Oz����o()�J���r������Ya�7��S�	_��r�� ����#�r��>c�B#vxd>{� ~��W}Cɸ9<�,x�wa�Ҷ��Ɵ'�|E�$ANU��Ӿ�PH�#lQֈ�3��P2b3�\�B+�Wй�n���M�=C{#ُ@A����Λ����g��vJ\63�!?LdP�f���	�;Q8��Xƽ��i�`\:���I�'.SlE��U���pZ6)�2vX��S��g�����Jw������Q-�vL�i��l��~?�Y����!>;�X���m�dwW<S�_�1 ��>\�*N�]�2hR�zc�u���k�l�V�����y�U~�οt؛���*�п^���zkk+��O��Vφ�c���zg�_Vhv���N}�38����WI M!{����Zf�-�ѹ���g@ �����`�������x�Օ�3��p0}~���p�((̩�]���a�&S��D��� W���J��I�����I�������jkjj�|�W�ؒ�h�LQթ
t�,��F�����j����j�a��m��1!�����[�ħ��A�?����K�I�:)�8n?qڝR*ۨ��*֭}�U�-����ED�c%abB�m5j��TY�/UA�yޑ��݁���bMUU5��M��Mu�@�Ծ
|Բ�[���dK��TW[/F@g�Je��M1��XU��И�JH�AX���H����6��hW�T�']���Yh�����i�(ѡ���___�u?c*,,�,�
��Μ��1{���a:�QWW'��,O��Դݨ�e�HFV�C:�4	Q�sVΟ�ι@{_�nn<����ot���X��.�Kgw�����Ҋ�g���R۶F�X7O�������`����y=.l��Y��؝�f``6����A���~~!�n��������6�����Uk�CMG�P:I
�
TTT�ݩr��v�����䐩)M���`�������խ��Ç�5��wNH��(�ԡ����RRH+++��oTU?�vG|������3�x
�?�>����t(m��\xo�����`��t���J\�H�.4�{]1_mf7U5�n(�B�Ǽ����������@$�����8�} ks� �!�y+��C�b�z��!i---3k��!��q��^��'=%���&�������k{{{[�L��.�5���	���~0�3¿��˨#��, ����.��(#!��O�mU$=m��F��~+�V88�[.}����nД�.�����=	�O�� j��f�k'h"�h��b��������N�4h�����!D����_vn�&�[��H����_[�o8V r�4ӂ� 
����ȱY/4dtG��v��6pۢ_Ͻi�ےЪv=!crq���zA�X�깙���t;�¡C�C<�ψf��������7Npf�=:� �D;��҆=..���III!ݺ, u?]o\=��F�k�������Ф#H
�]!�)�^)*�CX�j�P`��c��3`�ПB�wP;��ߜ�:����r��r�
���@�~$P�� �e44��l9@��{]�.R��u�~�ϖ�4:\��mq(�{{��b�uSk(k���z���u�T��E^}�ǣ?���eMW����А�� ćGB!�����;�K�o
�9�\�X= HIWx�;U�Ș�u��A������`y�����%����kh��X��J�ƠD���9�r��~w�K�=�NDӅ=�o1��*�	>��N���~�%|�=θd|�e�:��|�^1u��?(yx�����=%�HM�7?����W�&������Zr�3y-�����7�Ⱦ>~y������N�m����=��1��ԁ����׍Km�˲�ɤ�N��ɞ��Gp� �^�C4���Ϗ�yin�7���XU���g����A�]�R�Q����r�z�?�����,D�-,*Un���ȗ��h|�}/�M!��7��3��ƻ����I\ޱa��sZ
��>f�%�9�nz��vٯ�xHK�d���ݭx�ܫׯ�4���7�#��N�B�p��iÈ�P�������mY�A`���{
��s�{,�bp���X��m���җB����D ο8[ö����@&y���b:�QL��f�����O�OE�E��	 K`��C�m`��H_�W[����	��)9�6|���T�w���KB[;Y�_���q' ���/��a��b�Ωg�(�h<_MNNvk����#�S�u����F�"���0�)���!H�}c+��w|�w�ॶ���r�s���F/������0h�l�A�RY2����~���L����b*��v���B=��;%x%�U�%~�L��ODnObI���f׻�Ջ�,���aeSMk1r���|(��vw�`z�Njԑ�N��;��	���$"^���@��Ŧh��-o�{c^^Y�vE��B*u-��o��4wt��y_:�\x] U!]B�1�|2'
�9��-)
�TX��z�N]� z&�����XYX����_���]s�x��l���Q���V Ւ)�$���3$>xr��+"3G�Ż����E`�a��M�v^W' r?�UR�X� �:�)�ZGZP2��\.q�&_D��!� �$3'�������ԥm?s�3���K��)�.�ybϯ#����Y��_ ��5%����� ���Z��;$& ��->j���SS����=�;�N]Y�� P�g���`��v�$C���;	�,Jk����Y�2Y���N)��_/`���ttH�>:�4����!a�臇�����Q\�q��4e�C�9v���dr;٤�����U���r=�����{� ��Vǵ�P����^~aaL�o���H^@2�vm��~Cw�����,PCq�C@�ӥ�<dT/>p�'���n�T0���G�����Q1$\���k����}�Xl�L|!��p&�T���Ƨh���;���m?w�]�[ޫ^�ʒ]�x���K���X�bm�:�𰛼[K������/���@�`~���|Ϥ�=FW$9+]�ӧOA����^:�2x�πP�\�;㹬1�9�-w8���i�7��w{Z�ݙ꼠�a�"��b����&�۫e�����Ь ��G֍�	)�_�io��4��2Q�wA3+��}���'߁׭��yř�@|_TJJ���??�C�C�� �A���}ll,�Qr���*��L���Lsu��2��9J[�n'f�XL��K<��f2����w6ߝ�v6%'�X�`eł��2��7) � D���-ѩ�6��|Y����(��p���g�		+K�~k����w!.���lt��<R�yu�����\����g�;#�4ʺ��XS����J��9�u�/N����묁�,$�eci�9��p-Q;$�5v@��W��P2�3Y�M)Hi�E��DG]]��C���a'�x���m~@|���*P�??��:���RVQ�r����;P>�wZ�s��~`�<JE��?�;޺�J��j��t��ˏ��}����gA!�s���?���`
_�Q#�8@�E�@x�_-��u�
8ɧI/�c��u�)&�Od=�[HohL��hh �SL��%r�	>hv�X������t�a�����Z{SW��B���A��*�j���'���{V[�#�������}�,~/e}| ���)��҃t��ׁ H��)����گ߂�D�8�ƅ���@I	��k�(�yG!@Q�W�<���H�����QE��zX��.#3sg������)��b��������z���0���\�ҡ���ݲY��R���!�v��B޸�-H�k�����&�@L]���X��A���X���٬��G�~Y����}��r��~Ҝ��:�|Vc�?K=�a����MO�{�Hs�s���-��e_$ـ�����b��эU�d�ڗl���nعVw��{����S� e�̪X�' !s�BU��~.��cݨ6Bs�O���l	�i*�>kU�LY� ���7Jۻ=kob��7_L~}a_`y����|��;e%�<C"�%#flo�>�5{=k��p�6��.x�հ6�	 ���7���c��^���ϧ�6y��Oo��~������?��܆u!�Z��c��!,��]a�I)=��u�·6j@o7�gM�����7��u�-���d�Ѫ2Wk�͜(3�Rz��q�e#�ŋQ��p!,�n�1:��	U R�_�PˆL<(!�]��=�`���IC�u�e�!��ӂ;�1kCm�U��	�8Z�k~�ay���.Զ�Pȭ�H��3�����p�_��>�n�E����H�Sݬ'�F�~<[m���}������1�8e����s*խU�N9x��<����{�#b����ﾥM�����a ��*o�xIB�&fr��߿�Usu���,M}-� �� 0f�,�)�P3x!��¤ �M[>3�n�d-��dR\�
W�n������L�&]�>��Od֡�����p��4t�q�~1v�V3hж7������"C�r��ߛ������?O~����´&��� �$y/���]K����,L.����s�9�$l�-z�0�	{KX�^��!(�ZVx��j�3VQX���3Ὣ���o��e�?~)r�8�o��ihh���n�~ۺb�ANI�۫� ;�a�ӆ.����b	��v` 1 (A�����,�s �4�
�u#�y������ KnPܑ哪m��ȩ3oL����7��Ƌ4�{�G�:hu}_�f�8���h2@���~���p���V�g����0�O[�O��j%<��Ѱzp�H��]/Μ��<��B�{�Q9=-.�h���� σ�B/�G1~���&K��"��ݸf�,����^m¥��y�tnA.A#��3��6ףw?�%0�N�Ư����/�����r�m���V�}w�C� �yll��X�dw��5k�a�	�7���ȷ��bcb���222ڂ`���yR�Np��j���8��=�)�G�q2"��4!**�ٴt\�*t��`mz�Hf���8���}��<ȍ�.	������ ؘP��J|7l}�;UN�U�R��[Qm��=����ٴ��Od/��\v˻����BpN ��m�~{�Ր�h�s��������G�@��/�:	 T����~�+��봥:�(��G��y2���ɦd���H�6�(ğl�;�dde����h�?j=Xn�C��4��q�<3�;Ád.;_�q5����z�!�tf�H�+z�>��edD�:�[����!�L�u˅?d5���[v~�k�M7l�@4�ᵵ���gb����CHY*)�CT��1C�U��]h7�O<eQ%'vx=Éb-��p��>���r�n#Py�l�L�>��<W6a���&����5�UoF��r\#[�ed����W�|����¥S�'nlY�����r���g^��U-
_�DG�H_�y�t�H*o'>�Й3�޴������6Uc�-�$DC#9Җ7��g�M�L��r��¢���K�!ǽ�*�8棴H��q�{=��ͧ�A��H�׶\��&��;1B�����zƮZjj� 9Μٟ�V��I�Cs��9̺;:�f,���D��^�o4`�q��XSƀ��I5��c/X	���Y�L'^��U���Oi����*{>�p����+�u��E��7-�2�JN�U�f7��yB����W�jP/� à`�ffv�\��������J�Z��L��o�(��{a�m՞�"�s1�OA�����}8��({%���w O��@��[ѐ��d�<r�8ܨM��Os?�x�]��~�q�2z���(GP�I��)`tq�K���	��HNndc>sYLm��ѳ���t3��\CY��J�K��=��"�oF�'��B7Ny���n������r�G���c��EHj��{LW׊�b �O�W�"A���}VՓC;O$��0X�2y���C����v��J����+LWk7� �d�k�F	t�ҏPЅͪ�+��1�$.T�@���::j<��6�i�9���*L�jlW�&��Z}4�]��&R�R��86u����r��G���Ж������{��Ⱦ��%��?�6����1����)��� MW__�w�y�ZJC�����6ܚ�ӎ��C���c�E �D\J* �G�~����W��K�j�j�����+�?����h ��n�v�ٻy���
G�@��E#���R�p�:u�����xv��ϑ��\V6X0���}��Lܘ��Y�r���{�A$�=B�eƓc9t��R��E�E�+���Q
�A�a��-�o
.MQ��.ˈwW;_xm)��o�:? /��=���[��>8?�߅Z��T�^Y�ۂ�V������/�>��*h��`b�4��W�M��緂�x{T���9q������P�I��t��JD���ҔXa���_�������-�`t����xh=�`{ņ�|J}HH�NU��ٳ��R��kHzWv�'���y|�6��Y��?V��ą_�ѧ�wʿ4��Us e=�Y%g�]��|A�yu��-O�25o'�����C��?]!}��="��[��e(�fD���Ff,��(�9,��g�<��{ngo����3��)mk��w�E��z�|� ��ɅI ͖��/K�S$����==�4$�D8�������wHs�J��
!:��Vݵ�\<9q�UÇ��w�A�͐19>>�NL$��q��ӫs���{7�tz�`��AC�D~H����q�+�_��>92Rmm w���8�����L��L����xjY�$h.MN^�D��\к����
��TR�A�v�gI˟6�_9"Vw'8�I*����Yڎ'�K�!��\�o9s6���!�a�:��#��(�[�L�`�Z����#\ 7��S�����x�vɰ������<6A�&3�������
`d��!C6zu�g�u��M)�Y�P�e,�H��<5>~|8j�a�k2���л�Nh�&���gb$E}h��B^��ص�<c�����&��d�o㷒|��å����"$�+�r�8��w���h7x�	պ��D��1�}����u�A�lϳX*��M::�,�+R�˅�.0���k�~�0����ھ}�v>�_��|�<��@(�6�^ؒ��Q�ˢ��M��P�vRR��YW8���ck�tq�hu�fy�º��W8���J�W��֓�杕[O;`o�"��$c�-��Y�)��C�l�ѻ�CC���
��\��O`�_��~+m1r�n��������u�WFGG��8BCC=#� "@�@��7�g�_��'	|��g���N���<������~2�G�^���H�^��ȵ����%�y���s�H=�ٜ�؞)S*���9�jCb��D�.�<����^I�����S~E����s�+֩��K��u�~w�
��z���Y x|n.C����8����N{�O��o�آH񋛂����}�F)}����uI�m��dLL��J.�O�F�˙(� �S4B�J�Zq����N��`:H"�N�-ۥ��)JJ"@���q���*��$�e��x���8[Y�l}mm	T����o`�aa�?Ͽx�6���1�jt�\��Ŭ��EQ�G�+�
?6"������Ȍ��_��z����B��*y
�t�+*��Fi;�k@�wY��7���aPd���7P��h����f��׳�[y�����o�^� 2�ű��t�LD`s��4hg���~<��*| yD���\�b��\`y]�.7 xEꍥc�5./P��T��,6З���	�o����`9*mg���Q���RFL.{�)
t���O&,�>Tl�Z��)(S�S,C.��W��6b�7B#��N{m�8��S*}�>="k�����Kp���KuG��u��z��&S���=z�p��u�QRy���A3���JG0�3<�-�45-m���~�埯Й��Թ���J��[wװ��@21������Z�@kAs� �SDJC$����U�Τ�@�bo��ۛ/�+I�~��&O�4������ŸjP{�J��"��I�`d��y�9�_����䁺I� v����Eoh�������� P����%��"j�I=�A`��>$����^��	p2	�#L�_o�@��DP�ό�o���]�U-���qicQ�C�慆�����G8��,}z�$�j�;�;��+:X���{ 7'��`���b9���
e���9�g�>[:R�ի��Uh�Gȝ��B�s#�a�;pVl�c���� B!kі�Æ���H溆F*�^��Do��܅I��Eo4������	�*uX���^х�i���~=l%B`?��u2'
PG�7�QWţ��{�)���ح!C�w���d�%�@�s S˺]fV��Z,���HiM}}Wj��4l^������H����N<z/��c]k����`\�'zj�V�ß�����d�K��/����"sE��YdX���`�6%C��'0��{�J.hLJ�V(P��t�z�19���B�8P�x%9U����"�a�"9;0h�##.Իh�,6d�Q�u6����~�]h��&h��x zt,z�HЬU=F���N��Ӑ�msHBSL�� AOqa���===}�X<��f�G��%-��rϫ�}?>4���1a��/ؤX���M�˘8֎����gOx��.h8��6�)��p5H;ɸ�AI�r@y�΋�Yf74�g�?F��������}:w\�y}v�op����U#h�A����;Ō��窪�/c��ih.�`����'�!�f�Y�����H�!�;�$���p�e�W;e�{N� <Éа%�u��������U5�lB��Yx�_�n�=㞶:6��'������9ҽ�hˁ����W�h���oh��5��ZY���A��L�^3��p��y�Z��=C��!����M_y	*�\�s���@��O��KW��=�r�`�r9�p�z^7��^����s�,�@5Ή�X-mC�]]i3 ��.bktM����[ ��4���'������=I�FaPpiu���lku�pY�/x����*lĦL�*�x^�|�h�<�.(.Fw�w���Y���oR�xb�)\�� �Յ8��ڨ�N�T������B�+x��J�FLL4�0������a�.��ް�&U�|���3��B
�rL�d�LFM��t]��>�O#��ߌ��`�7��
`#���m������m�y��`:�֩(r�Ʊc������ s�SRv���h6��+�҇h�!�	�r��P+Rِ������)�v�ޏg��I��fD�8�%��f�?K�h*�Z͇$껡(
��w�������it(�=�n�R�;��� O�6�&I&������GF �f#�U�x��Z�Vߨn�n�[�LӢ��gb M�/3���;!0�7���� �[V%�$�126�=���]h�y�Kqo
kjϪ�-��mJ������(��X)L�,��ɸx�˸D,a8-� ��|qcF�!���X~y��n��B<�C���@M��Z�s�O�׳id��y��LV104-�1A`"�������t{��:�4�5JRBJ*K��֘Y��m�`$�^''��ʊ���H"�M������}����J5J~~"�ڍ����j���)��%��N�tt����x-���;�e�����R��_�j��p����%�a���W6B��������r�9���u-��(SM���G�ű�]�7����f�74�u��H:�\��"_��[�bvޝ:�}9;C��I��`ye��n���������H��/� д����f�������@�C�<w�KIII�ڊ�D�!��AL) @lkk������7P���- ��`<b�k�i��#��(nj���A��P秥( b;S�t���((��~��=2l��>�EBAA�qp� Lbp5�(r����0�w��/�@+�@T�U�i��j?~�xLF�)  Ǥu�[l�ܛ�6��8,�`�<���as��:�  TZ�����h3K؈qw�P�:���~�V��>W y���F�U$hG gg�8f�����uT1q���G�Z<�ee�~�ࠣ�?~�ʵwv">}�4(<ܳ��HT�BU^>>
!!Rvvvց�?�N���u�Q��@������cs���i\�������������TFN�1N[{��9�d�<Y����|ҋ���R�' �.�Z������p��^��H��Q���甊���vp:C��c�������Q����PˊII!�	�}��pYNZ��N���N�������l��b<gt
1��W�E�ДA�ƻxɷ����_�1QPz�p�5�/./3A1]n.�A��d�P6J���H��?WVVΘ�I�@��.P�]Z_G�-B�y.���e�Q��,qZZ�����27\��1���5�����[�my�������G����6ɡR٢�@���kC�.D��֪�Au��7�]�@�cPAj�=��B��y���𥡡aG��;�K<h_��%%""�:��O�q����p���7��ǗN>h�E��� �!n�5GC�\�}�`����x�������
:��_odN���y��QmF`	M�V���J�q������x�o�I)���wi�y��t43p�:���w���%t�刪��Z\XX�������W.��AH56
�������3��|��q?/���w�'��>5%�i�G��2�������x��򟅎�5�.t�z��w����:F�~��K�_����BPЫ8�O��
3tk����zch���1��Ջ	�]�A�����`{����E)(�������`8�BUaaa�6���HHI���"~��L�zw{]�#m�څA��$�W�L@@0V�GϨ � �xe�B ��R?�--##��HX��{bǇ�/��xgu����'&�-//? ���{
**x�Y.Gk(1��ؤ����K���\d� �@3b��-T-�5HΔ����(#{�����`K81�7���ڢ�P'��@־�O�ߥ���OMMM��&&&�d�-m@<cc�9��ˀ#@�_��=��������ݵD���h36!aPK�K =dT@�N�굃��<����g��>2#���
�������>�6B����G�n'���C��3�@:[*� ���l�|�"|�Ua!�dV�_��*y�����@�s655���>{�.|s ~����4��ح������h�	t�Z7��������9�es��I�}cS�G���c�jh�|����B��B+�� ���떟E�Zɷ�D�ں׷PCiB#M���~���Օ���&@tV��Q-�'vYh�孭�ͩH2��R�zh�sh����ښ��z�͙*�dk+eQ�ǲ1v䂷g��ຏ(R�ځ�Pʒ~h�1�	J�z�Q$`}�٬�~�B�2��x��a��a�b����#��&=A�fo?)�DA/�nNPh�"�l8��s�D�'ؾ~~J�w���� rBe5�J�8v*L� �/����|�
��u�;[�~�C��(�D��-�B|���tEG4w�6�A���`tTԶ�h��W{3N"5�,4������;��z`Zh�!���ܽ1�
M�����cw?�̜�ϧ8�g�����q��	cb|� ,,��ZEo��^�aX	4�<�C\]B�kv�s �R�D��=[|�3>� <L(�%\4���E�V�2M�ৼ� ��W:����E~ZN�{����Y�
�Ѓzg���r2��I�
	���;pܠFO�!�DU/�~Si6"v�B�r�&�� ������m9@KB��0������}�MY��}������W(�n���G���|��_l$�Ǩ�-�MJQ���J|�Rzj*�ɯ/7�E���M%T9�x�� �f4~F���O��{d�	��ǔR�=Y����H6PU�V�BU�ȯf�E�FY�v�J��-��%���F-��Ғ �����f�Z��v�X�;(8 �L�I,��@��7�8o��E���eJUf)Q�:�A*\ π���!�w�R���6^��8�����h�C"?Hf4�j�ħ�;�X\�c�#LAc����w�6hc6�=3W�5���O-~�
z�,h�*pp�֋M�lV�MBg����Y��dI��R�y��ABv�υ��UV�D��j��a%�?h�������o?E�h����ss��|D���:y{�(�h]v̏�����U������^
���ç{[�Jd)Q斐$�DY����D�^�55��	�`qkH���W��o2}���ym۞�A�f:�y�����Z?�e1�z*l�x6c������95d|d���(&&�n J�7𺾀s���؆7�h �*����R�4�9�|S��&�J�m�O�S~N4x��^�"��i���rk���٣��w \.����6KLF&�h��@.���`�Z�q�Q��{]n7��)�:��|��B){d*[ff�H��){��GB�
�PVċ��J�#{o"#;������w]]�K��<�s����s�s�G�
m�舞ɚ����2]��*����Q�@���|kf��o��8ԥ�����?Փ�qOS_��|P��x��M�l->!�胞c���*.��ȁh���۟���I�Ľ�P��G����*x4)w��^�-::0QBdȬ@
�@hI�0`�������s@��Ǐ������]F�b|��dEJ��o�Ϙ��|��	q�����A��!p����|��U8��}R�D�~�U;�N+[/�v4�G���p���8Ώ��5}�_�'v7J���W|Ʊ��Q����9���>{����j��c�#���������mM ���ֵ����宨�B��;3�E����:��遱�:uJ
<I-�@B b��֦t��93�F���Y��״�w�j��	��'g��*04�^���;u�!j
�,R�Ƌ��e .JO������JOW�\��tͯ@$K�=<���h(u�}��|�:+Ϧ�{og��6*u-��^'��!5��>�2����7{a�s#���̜���c�y� ��xu��t#�܆L���>�k^5瞈V��B��@�*���=�a�Z����{��z8p���k�#��4�kx8�u/��{�v!���d�~�����ԕ�'�s9��Xb`��{?��Ս6%�{" �Q����H�ͫ�Hx̀,�ܙ*���$`(�E]c-�?��{���O5D�/l�RV��	bPcL����������T���52T�M7���f�T-wy���P>b�1ͭ\�Ut2ω[��N��=F49�տ��1R��Ą�ei(8A̵���j�k-t���7n�:}ZÙ�OH�����Y�8�w��~4 (����\��ı��.���\h�b��
���sQX�`������B���<*��A�Q��J]�ƫ�����Y������m��ZG�M�ϰܣ���y��C�����c %�^F��y�d�����`P��a<U�5s�5��V76�7(H��·��Ŭ�����fӯOq���R�6���A���9����) &�

��?~������Ky���N��ւ�#6U%���� ��u|KMi111Aջ,�/��w�R�!���r��ٶz0�;��h�K�������He~�-����W�A[kk����T�f�W5PTpl5��#v�n�"����L9_�UGW�z�:sF��oFW��1c�����ۇä&ˇ3Xu}hq�}���7�Z@s��E0���J	�S���w�(hTTzl�l��گo|��Ѫ#9����K����L�t���H�Ơ �`f&2�i� 8�j:Սq���l�o '-#����0N6�H��VM�����������{#�I$�^))�D0}R���Pf9V��R@z.�$rf��vgF�H�&
>��!+/?�S���'�ski{o���cibr��yN5^��n��cǎ	���M ���+F)�(|����͛7}��������w�{�vj�J����s]��&�"����}0�����=B�d(���V�:P&�rGr�
�~�8�̳�7�1�<�����f'1�?,��%t��BF�g�~T��?�Tp^�Q�������Sl��PQY)�F����Ɔ*��+,Zh��G聉k�%���(
�{TbD��޻q�آ��L^\����[�3���å�=�"��*lzN�-��f��=�;��5�*�(���"��lx���ȟA�`w��F�\��(z�A������R�U��d�]�S��L����kv��I�ţ>!�6�իu�3�V�L�{qsFb���`I���ESSf�g �k4��E����K���zx�"�#�:�����C��A#Ղ�ӈ�,��p�/(s�m-m�7��1h�t"w�l��:����!�N�dI
�α�^�0�
���&�y�~���a�M��k�^d>>>�X�"�V��b�<�}�HЙ� �O0��KkX��I���U�X��X�'���f%��Kщ�����n��a�X�BA�����E?�w���#�������Vﳕ_�����<�a�p@^�4���'\=7*Yo߹�DN���	ˆ�!Ckn �d�㳳������`��|߸���a=�����<bf��(�ES77��e��q�(倪RaA`������j��c����u�$��ssxL	I��X=���(�����yy{��×��P$Q�ox4�	*���-��3fQ����3U,������d�Ӊ0��*u��h��8�\N}�>X	��ZE��e N��¬QUՃ,1�M�`����&4R�\�����#H�g�lB�[[�����-�s�]~��޼IP���n��˂ّ���;�<���=m����1�:#۫��Lt�fB�L�._��������6�zAvEy���6�ĵ�O�l�k?L�ٍSx!,,Lk�Is,/&���Q@`u$�wry�~�K}Z��:k��K%��������o�y��.\�yn.O��2�B����8HUvs�] {'���voP����+�;�"��	��V�K�1䘦��s�?���j:k�P���
�`����TE����S������h���`�)gEEEu^��[�n�{��x~��3
΂0����W]��{ʻ�������b���v^����JRI@���xu֞���	�ɃmӤ��?5��7z����ݢC4?a.�����l �FKa�X�'�B��}���|gB�٥�0�J�e�n��h�1�wX��J&��r��A���V�TsO���1^^߽U|Я��`Ӻ��Ɠu������'{s���@p|};ؖF����`ݝ�1��b���BM^Q���s����p�TG��+��!�E�*��3�����Y��z�4�l\���I�*�ӻ�~o�m�	k)%�tn݌[��%���ŭշ�)�[t��>é{����@�(�FdcP����a)�w7�s{q�D#��r��Ll�l����\_���f���l�4��q�1�^� qP߆��_=�! FO�f*�����/ǀ%���bTЖ|ͪG)N���o���/�q�p�|*'hX����[��=?q22H¢���a��<ioo�ԇ�>Ǉ�7�V\M���}nFX������l��˫��MR?rj2ZZv�e�Qoma-�K���a<��$Hx�J����:� �����ݐp�p����)C�W4���uWO��>�8�b�C�~z����?O��M�$2M.ǌ/,px	xx���(7��Q�����k����Qg@�e��tgi?�i~s|�����{� �� }��h��1�[z�UzR����ە�����JQ½:��H�{[6��~���u��3�\���Ս����7�����":���=��?����?A��͛�����]$���tX��J7�o y�R���oF��]�g&���$�xpc}� �Ë�R�jq%�ϝew[H5 7���WU�Ǻ0zr*
����[�I��ِ��P�Ci] ���խ�zP��/�DE���t�����=�b(���m���n������8mii�������0���	��	�11�>}�:����\�(C�5�����'*���R���׈uu3�ͬ�8A2��OF_�R�9�n� �j�}�$դ�R��� 6H�
��ˁ�>'�=U�MJFK�ym���W+k/^��.�;�n�,�ȜN�-!~���|á*���w����ܕ|[A�|�����in���h&���$=�u�2����7��F����g�������$<7���4������Kv�0�����*Ի/������D�4p��bnG�<Q}��r�Q���L�����b�w/ʀ���PcN�	u���t���𾒙R�i%/'G��I-dk�-���'<�^���[�Ӆ6<�����Ⱦ2l���y�f��(�����$��,�Fnn%����Ӎ:�.\׷�N��T�.�ŋ�*�b9Q�)à�Lu|�ŁH�Kn�A���k�(�m���+`�H��׏Vz;L�@����_6�D�
�\_�c����V�J;�ͯ��zm;$���}2�I\6�rejB;!�u�)�4<X����C����U�����3�*��n/��Ь��KD��N�B* W�̙��� kb�Vd���[�)pso���LC}�����M�\�����binaaF:��\o�;�-��9[-�������V�x�*�0ם�Zu�װ_<��yΫ��t��,����W@`�EN���m��Lj�?��Y]�{s��,2���N��Z�y�w�g�m��8/��iue ,��XHǼ�{&������k�vT9��'�i,�LJǗ�zy�x.v�]��b�` �r���|8�,�p�U�ye��<�W���uZĴ炚h�/����$A���|/^�&L΢G�����;K��C�"~�5�a&�DX*��]�*� ����2�?�y�^�eWK a��RJ��+GV�v���ݛ++_*��=߾zEv�޽��q?>��؟���, ����'Љv$�Ƿ�v�G�y���43�������Z��{�}}�J�w7��c�FgdK�V��{s�a�ӯ�>A��ޒ��b%�n�Br��`r� ��p��j���3���
Ƹ����Դ��?�Ɇ��*�&~�fǒ�;v���g[}��Α}�g��'�:44�c@7��5o�W7Ԁ�����|�lc���a����.㯯�7�	 v{�>���6��&��ԋ)s�:]ǭ+�߿gD��*���̺L���B�>���*�qRT\B�^�"z��}������y�cHY�ꃚ��L��g�@3K���UB��1u�FaQQ�2�x٘�KK����$�V�Wt��h��	<x�(!L	J�WN��T֏����\��C��/�a��g�Jo���s�
�gZ���$m#.v�3�9��{ۙ�؄���D_�ێ��c�k��-៣�f:�F��[�@���>��J@���^%��|�ͨ���w:.���2.�]���#8�`8����=��r��ethF�^������&�b`x�hT��/��B[8���ƽ
7X�o�
�lgN����]]k�$Z�O��F������C��t�墖�&E��P�亵�+�2h�C��y��4*�����@�X�s�U�>?��[gnff���s``J���% �P���A�䂳(j��_d�uE�_mrQ�Al���;���/�q�: �O��%`͡;k���+�8�]��epP;�@��~J(�s-�����$�e��d��kkix|j*��r-e�(�5��U��.�6��FP�ȶ*�e�o�D�����g�Ը������LLLh���ȅ"1�8\N�2!�����)��V'jQ�5�?�G}��΄cuQЦ�r�}l���sxhu����&��o��ډ�l��+����ܢĔ{��'�;�x�s��+�&+�b��Q�ɯ�W	�#C9���B@6��
�^��� 
��"ex�?';R(H�=��y!T�{�ޠj�D��ܹ' HP;8`c��[y, ��T��:NX���xu�B
�^����8�W�b`�.�<8��\�L��R����Vَ��v����ܬ�˿p�/��}5�:�nFK�2�h~�Ɉq�|��÷�ҥ7zI��CB��NS__*��c#�j⩾��$�v�=7xhr���-���[��� ح�d"`.q��& ��/aDDD�|jc�=Q;<L��-�uӭZ�����s� W:��x������dAB��"/�5.��i�-!�AXEI��=I��򈄦��l��j���f]kS��A��ĩ��[����Z�Vs�jiN�i�~�5�6(�t���)p%�D'u2������9*�q���C9�|�&����������9,7����3��bLxQ!����	��R#$�2Ɇ!+S��3�L�K:r�5'o�)޹s��Y�{]�U��m�������]�rEXX��%ע%�xw�7��u�J���--g���kr���B�}�PK	�,�]�.�~�}_���M����x��y���̺���By��"�����{;k vv~y��x�۫��m������/x�ֳ��W=��]l��y!�;X��E7��0��'
�w��!U; ����K4�r�������Hh9������І�q��G_�	�ڙ~-.�x���$�Ã �o���W薪?������ޞ�ǻ�~fi�}��'������k�22h�DJo�疚؉{�,wb�{~�QL��X���Y��l5�*))ͷ��	���v��N�����4���s(�K@�+�z![��}>����E&�~���甽YmB��["����F{;0�Ӻ>�ס�Q��T@���EW{��	\)(��Gqh3˽P}�X���'@�d5�ƒ.�?��ZBQjϡ��F���8�����㓓���Ƚ���o�cOA��Tꕨ�Xm�6������>�Ф��m﻽r%����o�i�	d�q��Ly��!S�%�9�����nyT����bj6=w�&�޷�.�9��PDGF2�kW�=�7%S�c	¢�h���x�T�JBj��{�4�ؓ���P=%g
:HK?���5j��A��ƍ:U^���}||�����i�������V�wͽ)ʹ���jҽ�}�j�>���#���ͷs�����\���8�4X] Qp��GƆ]G)hU>���W6�A��_,�/��盃Ĕ@'= �	%k����W#��w��s����技H}^)X��w�
�I}\�e~u[�Mk~���@�N��5�ٵƋ���m�~�ҳq?��<����cȬ��C@�n��n0�X��&6��ߣy^;�I�(�٣7{~ms�>E��]�0
�` ��mNʣ���[�>�d9����奥�*Ln�u|�3��U��f��1�'�L|�fc��,ٲ-����[��,�X�z(R��n~��y�n�~�4�����w���s#�媶����P� � �߿���-gD>���9w�<Ǟ����ם*_ �Itn{�{wq�h�/�2�f5�͢5>m�I�Pz����-( ���G�����d��$�Ӻ�*YX\F���)����` WY�ѱ&�c�f�����H+`�Q��"
�����T���Z��dԲ��tc�6���5f�R��R2���K���?X$�z� ̫v%�5 �5\�r�S�c�������������|}R�?��LF�ڼ� A�슲,4
�H�{fA���R����E��{N�`����y��dy���A�v��0��0�U�����0n+c~^��5��\�(�C,ԃ]�� E���A�s�EE�V�Ͼ(x��Q|J
31]���fƉ/
�-���QRyy��(��sq^-����u�*�	^�ՙFĮ����h���"��%������\��'��
����v��D!�ΐ���Ab�t����)���j��|�?Ѩ;�22����/6��w'N�ǌ�)V.>���E�5�9DY@ړn�PJ�Շѓ�� �����r]��^�{���3�D����ʭ�������^^.�3YڹB��t�׵\����efzKIK�ih��ғ���5�������o ��Kt��.�j�>��*"ҟ��&����8\�2Q�<��TG���:x\�c^(�onC�����)�I�n�P`��|�J�*�v=J
-�����`!3]����Xդ��P���[{r	Qu��rRܿh�{sQЉgT���@�w�� ���Og�zr��tD�s�={�{]]��$�2��/ �x��r���^Ӌ�ҁ����[�^���SR��o��X�de=��ڊ�h�4o$֣�#��4������\n�Ln����{U^�Z^��!�~9Vf-����M�qv���-9.ɾ[�+����$����_`�/YP�:�utt�t���)��ѻ��Q_Aoi���.��{zx$�ɱ���P���>U��Y�q��r]���故8P�m���!7!��2;����W��(˨��qrur"è��:�(�y��D��^�u7�L����؉���{c��Ԕ��7��:���>�ڍe ���eb~�d�͌�q���bk�3M�N�mt�-��[l�������7�~|�8�ڈ�L���̐?�x´A�I���'�o��R�2a-е���H��N4�	��}���B� �5���'E�Z5���5���8�TQe�ˍz�p��$���d�*,�U��F������b_G�V唎�ڹ��+�!�wQ; 2�Խ M�a��i�i�(d�'�(Cy0��2�s��Ć���B�é�6�����*}�p�K�F�g�!����]��lX��Vo�}����z��Ȕ�I��8��n�4W~���X��=#J{I�C����z3���E��$�x�Ǯ(ǟ�V���F��1����U�G��Vw��D0��>�5R+���[߆�(�]^慔���d+�l��-�-��/b$�ʝf�7�StD|�g�����s�����i4?k���gR�g�,a�L�{�[w�6�U���hN@/3����b��z}jT�o7\֥	���4���Bu
yQ��N�������^[�4��d�Jr��t�A�h�f:`�ާ�E5z%%�Aw�O��e�\h~���S�QN�������
��n����Q�n�?IS|'��@�;����j�#sm�q%YZ~i�YJJ��7/K�=<�3���꡾z5��]]]��Y��{��O���I����FA	uk���.��"&���߮�ޝ�'Oƒ�X��@OO�Z:b��[�vE��d�(��M���=W~w�agǻ��\����F5:$�d�$�������������5y��j�w�3�����٥k+*)��ѡ�����������O�W
�ţ��UT�;C%�����Tp���֚��$åo���D����D��2@%��aCx�֕}Lk6���ff��[ܨB0����n��w�a�!<5x��ۇ#��=�ߕ"v�U*="���+�y��j��h�������a��XA%�P��b�@�h�����e��TTϱXN�E�4S+���'=/6(ϴ��'���7��̹��J��l�b; {�����itc^�z�-h�VS�.ڊ*��J ?f��V��2=�2���یٛ����!$�*D;Α��~�z�����t�K�3`n#�� ��.���H���`r0HTΐ�Wp��oް-�����@eil�M��I�_��ܳ��^�3J9?񃍻{��~�O��5�����A�C�͜�DO�sHՒ:J�,u�v��{t��E6:��9�����e"�h�2�[�?!����ۛ�!�w|]��!R0G��q��l� �F��wI�l��h-ێ��k�w�ͳG�wꢉF���;�=������QA�[0<D��+�4j1d�K�))���t�KJ<o%<�����BЉ�ث��I�;o��g�bZ���x�H�,5�l�����9��/���^�x�������$�l2D�;u�E<��L%@ֵ`�Qh%@��u�>x�@��D F7b@��"���s�N{̶&��8J��%����5���A��	���h��gZ�Z
Z��fo$���!]F� ���x�&�$$$�.��02��2�8.�p�r(�2�II�	b���S$I}�YZ%�����p��Xď�B�(ɫA� ���p��aYk��ژ��E�沋?�O��H领��z����1bY���Q"&?����ئ���/!J�W���?�2B��Ҫ:C=]����,*�qК@;~�HC�gOغ7�k�/hT}ី�ų/�C�~� ����x��"��莜jZ���xݠ�=���T��-AZ�K�Wdd�jkkq�_qW�켼(s�m��
w~T17e���Pж�09�Q�H�w��g�������G�5?ED��yg ��Gu|�������ݍ_ݘ����Qn����%���X$A����O[�Q|�HD���f�ho��4���,p��ɹ_��Wh]joߛC�}�䂸2 �Z��㤾ϟ���PRR�c��r	O�Tڎ����6�9;u�iio�7N UY��zLz�kg�9
�PZ�����i]궶�ۓ��'E]O]��>;�ê���� zz�}��߃�Q�؀��I�����`�«��V�њ��.w�����O��'p�v�L����.��R�Y��i�O��h��M���:#����O~_�����bk��tf�5aDg^�:T����j�(�T�hOȶ�	���(�Tz�5�3;3o�~~��`�+��%�'_�i�<X�vY����n�F��W�E�j��nmV�@pH(n����޲�b���p���)eo��O�o��2�M���q�k�6�ƅ؎
i�Hph猁�
�ak�m7����ɓ脀Uߧ�@�t�<��2��[��5���R�5�@�Zd�ps�J����CL����P]-��=;s�M�U�Ë������l����]�$��e{8���p9"?~�@�"-#�4�T=�6ŝ���pe���(}0��2CCY���e	����ĕ�5))�Lͬg�Ba�;C��}oo�}�ы�yg�ֲ�M�1ų}e���r��L�;�j&CZ�+FjLi�4���S�F<`Q�ݮI~�Z4�4b��ӓ�Z�xb+y7V�LЦ�kޛ���֝;,譯�W����SGG��qt`��I��7$�i\�f��~�th�:�Ą)??ߑ�Eji9����9����&����e��&���z
�8󊋨rb����C��y-�)���4K�5r��[��] �+�n]��쬱��gՑ||<00�"a��ʸ̸�Y:F+�0ne�3��L�9�չ^��:y!b;Vq��q*��.2�i[fݜ��N��Ao#B�(l�հ�bqA\B�e`G��e�o�Ψ�]y�~��qbb�=]�u�Ѫ�A�s��g�}�����S���O�Z���ܡ����'�a������9�H0���S	�1��Ȇ(?��Dr�K�(7���l��$Mu|P�š���H�&��Qc�������Z������ʡX��o�>9`��M�%�����ը�|�3���d:�曙��N����9n'Ev]h�K~t|��U������� ����+î����P�"���C�5gDvq��Vz�r�?��}�ϧsY�MPf�����+����M�\Jiv(C���d�,�A�{}�iw��-�bgv�o�P�S�ӗΏ�h�=M�A]O�mǣ��A�Ol�!�"��gϘ��;�O�ͱ*��[;e�z�~Vժ�-OOZ���:�fM�k�C���B����Bd���E*&RR thg��j�2%�^�`_�@���|��~�� �t�
�>��h���S�r��c�����g�>�dA;Hω���n �EDu�Ү��c�1�륻�
cJ������sfO�F(p+D�L;�O�eQ��G��N�Kց��No�ˣ>��#t�,B��>չӋA�$�yx�%��{��0���=�Ø]=���%}�iҕPS�6ԇ3��s2����S�_>ʇ3�������L��7����0�]�p�fx��0���}�/s�u�X����H�tď�a��J�1Q]��X_w>��G�;�9'j�r��uv�
T�>ב�W�t��a���Ǐ���"T�ٜI�uH�=@�UA�R / n�ڥܖ�ٶF �a@~���V�}���\��n'5x� ����ꞁ��42�����Q���"��[������v���5}8���`��Wy�BQ��{I�*��+P!�`�/^�Nz�����r^^�tu��3��g��"8�")�Lr���5���b7J��������n@,��^�Q�ݩ~x��4�An��wC���F�֙��h���o�}iy{���s:I:0��9��T���[��Zw��|U��EϤ_l7(]�0�������DV�L,���F^NΠ�V��P������c��߃28@,5�p�8N7~�!�����9���l���TEg��P���9����5���2RQQ���###�h��Nmm���o--\�R��s$�������w��'�J/�hrJ|HVJ�BwD=����)��|` &&�T\,���Ͽ�`a���S"/L��J)YYj��K
w�.[>(�n����-���e#���.���)��q��Z
�Й���V��K
�8��F� �e�H���������=&�ϲw���fQP��
�l��D��%�P���~_C�Y��2�~\C�R�_����a�~��å��}��'\e��Bc���š�c���z�ݤi�2�i,�8=��v,��k˘XsvӎK���xR0s��b��V����G�F������3)g7�ĉ�==w�q"5��}|N��J�揇|"�����"����)���ٳ���b������Gq�4�^��a�#���R��N�q	QQQ�/r�w����!���3�}�ɰ ^���������sa��>8O/0��d6��E�H�<��sl�r�et� �P���9e����
f�H�1�и+F��7N͑�g �55�k��OR�8�Zbg�x�*��=�P����ۿ}��h-��a��/O�	S>G��V$�@�\J�߿pۿG5��>Ak0�3�HE镬@��(4�66��`>�Aб/�t/�@�jh���s�����Ԓ;�,6��;�DhTV�ƙ�2�?����ë�~T�r��u��?&��u�틯s��w�o�L�Q���G�3D��-�4�h%>uZ	�ُVy�d��,/����uM�K�7]�9z�@`e�×���X�;����=��#���	�D�^�Պ��� ��+7�9�Dsd%�.)F�D~��{*�"���S:*N\��wt�;1,
'`:�_xE�s��Y���g8W}dĎ����fb2yNz��.̕��6 l�����R�\V��4�T��z��D"����2�����dŶ�Q?��^B�f��F�u�I!��=�(6>����^�]�9�B��M��������1i��ʞ�*��`m?&�����p��������@�a �����u�iR�������8�M�B� ?8���E�k�OUU����K8t�4G�옏�5+���U������>f��:�y���g�S�{rݣҧX�΢�]#������[����.���H����,A/^T��xf�͐ş��ξ:�}䚲p{T���9C�n����*�s%�E�߇[�p��W��=�ϗʳ̓����g)F��O�����-��[���~�����U\|/��қg���њ���x�����	w�;jbuV���OJ�*�Jű���-fff]Q�/Bg�v+��e�H�R
��Gq2�n2��!��K�F�f�:�~��FG�KX�q^���{پ�U3p9y�+:�o�t��S@�UE�(�#��$����Q քl�r��WZ:T`4��D�535���v9p��H��B�g�//�צ����ς�Z�@�|I��))���U�M3�j\Ro��N�m�T��4W��W���q~�25�s��d{�	Fq�3!����{ɦ��b?��������DFr)�4>��?bkf���hC�fg{�E����X)t>����
��8{Ǎ&m�s�;�l���<�5�,%���B��X(��i���Żq�_�ҿ�ҪN��Y���F�ٮ����%��o���<Wr��	���@��f9F\�P����NԊ����Y�R23[���|��$������s>�W؊�+�y;ȐN�_J=�t��V��!�-k?o��ߴ{#���}�7���k�}7	+�Iܢ}r�s�]�7X�cq�j4�����j�	c2�Q��,�#m��� PK   Pn5[���8  8  /   images/864a21b5-9f7a-49ef-8d10-822baf4f1419.png8�ǉPNG

   IHDR   d   �   ����   	pHYs  �7  �7�݊   tEXtSoftware www.inkscape.org��<  7�IDATx��}x\յ�-˶�m�[�w0�@�`Z��J�M}_����r�K�/_^ 74��1l�\��ޫ$�Y���FS���9{t4:3�#��z�kΜs��g��W�kۉ�O�>d��B^����������<�����5�W���vM�͟B>�aYY��O?�L9[322�n�����}�ǭ~d|�ݏ �c|�}�w�.��ݻw�D=����]j�Oo~濥��<��^h���t��ijnn� �����'��{�Y��Z�Z��x��ɟa�x"��v�V�5z�ر�Ç�cǎѦ͛�ĉ���DWx<��l�	��g&�����فA���3�$QAX_�k��9��F���T^^N�ӻ+O�Y�t�ĉ�x�bZ�jEDD������ύ������5
31.�|�.@zz:eff^���uΙ3��n�Jn�;܏ �_��T���M� �!�xLw��&y�PF=��t�O|:�/���A�G;�u ����֬YC�!O�+N'���Q_`111��]��(��-cfTVV����7A��iӄH.\�i�wPv߾�}�_a��dH�D  ��t�) X����@L�Z^J����Ma���� �kL�.A��)%8K8����+�)A\n��Ϊ�˥��6�5hC�pR�@|�Fet�'�! Ѵ�B���D9�޻�^�W��v{�f8����F�L���z�uc�QB|4]����v����L s�����h�8q"EFF��3t�Pڼys�N�@,c����㔑��\�t5���iԨQt�����ᐾc��[�N��@DN{tO����Sj�8��n�{�P~A9̖�� �� !!�����F�d�=������c���G�N������ޔ��	���4b�_��n�=Z�|��>�ֻ����ٳŵr5}LJJ"�j@�[ll,��Ԙz�A��^�����M����b�:(=~�T^�L11�roQQ�F dҤ�t���>i �N;��9��S^�L���X9c��n�h���Sd�)��WFPD��Y2z�h�ٳ�Uc������@�q���kfNnS�t���֒�FEF�?�=}h�{��Q߾}eB�={VcY`7�d�xx��!�� ���z�j�FE:����tj*�!�����j(��j�����d!�8KKM�YG �4B��xiJR���"�ʳ���PN	A��@��8�.'EGE���^�~4?pHCC35��7'(\QQ!�5;X
�٫�.x'�n������E�N���������pig,��Ϻ�F*��%m��_~~��@����H�5}�����|�z�w2q��ޟ�w���y,F	:��{�	/T��-��"ǚ�e�~_��e׮]�p�B�nxW�َW��:92�n�.cM�]��&��6�����#�[�nҎ�,�&`�~�� }��޷GD�o��k�m�N�V`�]�c����Q2�������G��?1�b���jcYBx'�lp���v��ؘH?��m���03�1>7l>�WX�ܹ��ʍ���Uk�V4�6RUM��0����T�z��**NPU�����	���8K�d��
�2#z����{_.%%�PMm#����s�63>�m�k�PQGe�5��:���1

��l,c�>�_�1õ�+���3A��Z���Y\Z%�\H���)Ju�TV���J�	�B���J��Ѹ�6**�٢։�X����l�8ɉ�'�������O܍AЧw�Ne����vYjk��9WV͖;	NT��nǗ��41v�;Ƙq���Ҡ�=ev�u������{�/!���J�=��Z�җ(g|q����\*|�����1Z�6~�h�2<Uܛ�e��\��>+Zfgh~� �ҜY94nT_�v���cE��L���"I��ѣ��E���@�S���!I4|h�����������06���,G�~y�T�
�<��������ѰR9OfQ�Dʌ���WF)��&� �Naʱ
x�)�f�{̆�XF���w��Q}���o��K)77Wp%	!�|}}����=H���q/��(�&Z�vy�ɘ�iۉ��!e�^��� f��3�@f�ρOWl,���
a�Z�C�0#F�d�0��t��[m<���\���9C�o;p��ggӠ�E������Z<���"�(� ��Rv�º������(,E�z ��	��١�.���6���s�h9�=ᰳ��H�U�"K� *Ax�5��M��6��q���m��7�7�TP[�.eI��>��b@���%TUVRW�x0��"�S���fv5�G���X��}�0�78�G�X���-..�)E�m8Dߛ���L1��:�����G�+�L�})��oma��(�>/f^��0 �R�cd[�'��}yp�~��!����"�WRR�ɐ���S�^�$㼮���X��ƌ�cON��*cf4�U�����q���J 0:4������w�˲�9T��������Ί�lX�x3M�/�{��a��νZ<$66����'3D�!�nEK��Q��jZ�j.��wC�]E5��e5��+ڑ��U\M���	���6���^D�����U�r��N�U�Q��;_^M+V푾+O8����m,u���C�n5��́(���b�<��Ю���������'�`�������"�˭gb:.Z[3^����`W 8���k�6B�ٔM�/Ԋ_���"`7\��$��F�����p`���E��P"�Z�m�C؝���L��{j��řeQe5��=�TPtA�G�aYJgGVcz�Xz�I�]`np"+��p��c.�Jx^��.�xݭm�D�g;��g�47��S�"��ϢP�h���hu@�^=�$��B�Y	�a�3b��p;��˄�Z�\h�r[����TҼ;ǂ��65�o��q��;96&ⓙS'���Wԩ \�U��͐������,�G���Q�Cu,2"bbbiu����C@��&��^��j���FE:V̚6$}�G{hĈ����'�ܗu�09QB��@i��+�ǻ���=�AB�� �OY�fBZ�E��_��|�sj�?���j,�_Qyy膱
�"�g�:nb5i���-��R�b���ٓ8��k��P!�Ʈ�c�2QQ�ᚆ%�2��jh�(�o ��)��aMCքQr��G��=mf���7c[*)#x�H�QQ�L��B����YL֜�팥��5�s�e4z�x:���y{խ���h��4{z�M������lQ�͝�g^�n� ��3�X� k� �/��9ħ gZ�����vL��x/59m��2'�,5��=\ �p��a{������9v���G�;�P_/�D"�q#
���0�bs)E2o5,뮈�]�M�}�-��ɞюi/�¬�����H������#�8�35� ���Z�<�23�" 8��	�����;!�=\��(�
�,lE� �!RP


|�����q#')6&��v��&!��4E�g�!H����%w�Wd!<5�I��5m	�npO I�s�z+��G�	�ZKף�����TU��'O������1�����Zq�]j7䎓�q3!l�[k"	��<[�C+��؆��!J��1<8��^�_M�p�OD_�C�6�KƮ�;�5`����wV7J�C]��V]T�À�G6��C�Ls�<`T�?�3�� b�z����B�0
U�|�
���18� �Pf^^>��ӝ��ѐ�=�e`\�;x�V򔻔 SH�'��Ķ-��f����tO3��0��LY�QЖtXhάaHb��m����t�>�OH���l	JC~�e��3g�p9,���X����5�~U�6���G:]�R�\f
��q�QA/�����@ ����6i͘2F�'�g��n�q~�648���L�F�j���AD+=WD������G�sh�;�����ÇdNܲ�d�B������,=P!e�X�kUA�̣�<��i�b�!�ă��#Q!\�X��}n��NRI�޷�݆͜�so>����!�vͣ��N||��gU�na�֡;�u�Y~@��blOu�(��@NF��bVFe�KW?#T����ώyzU���Z��^�|�'�,a)\'��^�
I팤2����=����[�˷!�� KGB�@����iÆ2��!�r�ٞ@�;9%%h���$��5��*@���{� �Oi2-��L��⦦��v�=��m�1^G2�)��a;��mW�%�W=%���r#��XMvOL���Z�/]č�.�Pk]��H�^�A6<R����/�c4�մ���dB������B��@�J9	�M =++���0�f̘A�N���`��@�tfzJ|BB���m�Z,��P�0�\�[��ev-�D�����*zs�&;�ODRbl_Da� ��#�wtȟ:u�P��'���M�BB��X��B<��1P�����P���:e�,.:�l+����)�~�ܹv	�WЂw%�ɪ�*6����C8�m�kK»]��h�y*���b�J�bX��^\W!��7�"Sѽ@��`���+��#���C=��X��D�|'^w=�䓴v�Z	wwdp w��?�tw�E�*��x�Rz|�����6)�ti!\y��ki�9bQ#��~<��8��aol�h����Y��V�%�<!�SJf��J��*�u��!RZZ�a�X��9 �g1��z�VQ?�(�Ow	7"�.���N������O����ci���^��<�����6��Mn��;��?�DK��a]�y^�o��f'kyn����&_�蟓��a���+��7n��&M���N}$+u�#��ì�ՎA�B�&B����
+Cߣ��L�<�����y�L��������쓕�3h@��w�~Eg/�̺���rxx��ի��h�Zt��5k��.�#쮹�ΟX�H��'��6�c�k��8��m������'#d����ܹsE����'����0� ����:i$M�y+�9���x������9��|���#QB��I�.��{��߬�C2�}���+��	�%H�K%e��%�����7���=��������ب3�IZ����L ����E��K�,��lh1
-m���}<[�c�����֟��M�������;�'Qi�iɯ�V����goMM��It��Җ�Y۰� �.���t=�n����.::��g���%_	~�R J���0]�������b�׉���k��xWu<�6���`��Vr��%Zi��R(!P� 2��w~@�u�t�4����ޥ97�&W�9*<{Z� OS>Y<���c#wm����%�0���"�3-QB���'�(Qo��1B���/;K�6	�*K=))�g�M"\�Q9Z���e�_ !:3���SA��B�P ��L~9~���Ȩh:�[F˖���: �J���3�X�ă��ЁC��F���Q�;���9�a�PF����;��K6B��U5<;z�`�ռ��R��{8|����sss�w	��sV����=j���N�v6@�"����T:�.g���)&���||*��N�>�;��c'u��1�F�p ��s��Ȉ�%<��!�ۏ/�AocܗK^�Ϲ�,u.ް���"#hDN�}���n�[����nW |u���a9ݺͪ{5�Ly���t)�����8I�qQ4vd�{#�{1k�ȓv�G���mcW'|5��1�V��+gbc�.�T���vh,Xj��HK��`S����^}Iܞ={N6���1��O?ߧ�p� U�J��4���s�˂�|�Zu�,�uc�h�p�
��ױ�=}��%�V�c�z����10�M5������Q�6sx����*���O�<���҆0�p.+#E�YEU�x+CV�p�&����Ӛ�+录���/�y�y�,<U8��O~B_|����=O?���_}��6e�5刍��8J�R�3���p5�*/S<׎ƆB�Ѳ����e�.�94�=������|-�b�%A�c�,<��؎�����y��|7�̡	c��|�W�M�Hv���#Ml!����!�@�y7���#�@;��5�Y<0e�Qbcæ#W��e3^8ݨ�"��3���U�iִ������s8l7N�~�ޛ���A���Q-�L��t��[���4x@O�p��O��H{�����C3&@�wt���P5蕏-P��b�(��X�bu���w�9lt�����q�~ෳ����xL6$㖣�*ċѪfFDD$y=nb���\�h�S��:�	�cn����0< ����cı12�=�|T�w��ҡ���{�W����l��B�H�����ЉNGy�܂��p~�u�B~���d��������m�y\�C��\��Һ�*��<����7���b֯_/a����r�D���GB$#�;�馛�;F�Ҭ�7o�l>�x��%-!�j�7�g�&�|yr��ְ��y�1c��O�Q����v��M�6Vу�'�������x,VKߊ�:���GB]�rEf�믿NK�]$�`=�<��>�B�d�(b�sf��!܄���U���2��ٜ�a�Qf�_��e�Ӌ�,W��N��Л�7!182)1�?2�b��B�E��2s.��� �t�9�D�-���MS�/�[o@	2f�@�ͩЁ�3�o���&���-n��n�}Z�6`Y��|A0�������{H+��Cƌ����^*��k��Y�b��h]W)Z�ֿ����wAIX�+c�Bp�&��di4��>ޥ�pa��5��"�Ƣ���n�������W����FʩS'}nkc��j�<��3!P���1���Wf�������l���6ݰ�*�{����ҙ3g�O��iz�����
*���������ߕ��;�M�MI	1�*p,��nж23{��?��h	ΦF���N��g�:����IR��b9��R�я|���2�v��E_�h��g�[8�e(-zg���*�[��{��&�)l�#�7-5^�0�ڗǬ���LY�	�.u,���\)�$Xe.�j5̮N��5d��^��U����ZUE	m��_� Y�u�9�j�����!t�����}Ǘkv ���5��\'K��"Q��E)�U�P����aC��%�E	a��"`����5��7D�I�Ecƈ��H	�V�Ҁ�b����쐞={�������٦f׭܅����?�9uH�;K��}�$=�Ly����M�>]~�L��k�t ��Ŕ1���1G������w�ɣ�x&h���Jߠ�N�7$9 �����]Ͷӻ��t&F���z���13�I11�0ch�嫏H%&p�!h'��LLI��B�L�0�	�&��&���_
b����wl�O�հ�A�g�T@��ɢ�|�Okn=kE�F���7��/��\_�s�����\T�p{��.�(/�����Ԕ�璓�tW?�um�Cϔ�$&&r��S��k�nr�t+�u6��7��B�镚�z�-5eHo	@ ��N_{rQ�V��̇"��\D�Vیz����ȭ􊋎����Yz�=(�SN�}�G��:AC����y�X͘2d.�\��p�����&��Q���)� Nɧ:�NqA�� �ZG��ڋׄ�Q���)�	�K>�w�h�nO3�K?�ޖ�g��&է��*!\�.������76�}�����q�d1�i[UU)�����W��7l>&�l��̇�CMM.ڼ턬$5vOH�I�>.S����-��C-*�� �:m���d�Cw�-��G��n��M�'Ѹ�pDUN��/Ш�wRl\����^��*I�-����\7�o��ZP���8)[��{��a���¢�a��<�0L}�>�]�e-_�W����J�*���V&��x���g���I(X�?rfԽ�XGH-�./5��R@���V:[�(C���{Qm�����.��\-�k�f�:���+2�S�8�Gr�w��E~��6P!�`���R�+��"Oe��J���v�X��9�Z���׿��3/��}~��a4!�_|�W��"�R:�mJ�P����D�������-�Z����w���.�$����P�)�F�J#5_.0[��*�@)�h�ȗ�܀oP�TE�
���ǢO��֛FQ��t�"���yR���5����+O�
?����C%��b�6V��/rjР�bby��cY4��k׮�铲i쨾 ����ְ`��āw�1U��r�k��* ~'O@7���Y�Y��҈��۽�/>Q%j�R�R��2-�������
fa�6�9�X�"���9��!ܮ	�:�((
�A&έ�;���W_9,k�ރ��ֿ�}�p��B��wV&Y�U�>I�@�g���_�nׂV��'5bh���C��9ب n���\M&�TҜ��R��BE7����=�6�m���EB���6�j�x|��������Օs[�p�uK�����L��of�f%���Z&�V��0a����Ʌj�5�WLL��'�ۭ���U�vei[��`-�2Ly�፥K�U�'�Ҧ��	��
�����M���Z�ŏ�lv���K
L�v����m��7�����I�у��ˎ�g|��҄�2\����ť�u��=�"��Ӗ���*���6�|k��<�ljJ�D�X�U��sK�<
��e�?c���X���0�6��o��dMb0�n#G���?����
W�����eӜg�'���S�xC���q�t�N���p
�U�-��`��)��{7]�t�d���/u�*t�����ӟ�����?�vp0�S/Q��ݪ�r�zh�V���P�-�k�|@����E��O������u8H[jǷ�p�\#�dLς ��	�x�̙���7�v�4�GZ=��#t&7��n�ц���Pze8�&�!YY9U����c��|m�{Қ��k].�6�;j�b;A��sv?ڞ1m
�t�l
�h3''G�A�)XyS��s�}����WX8����I��ʦ��￡OW,�/7na��:<6%9�*��)..���������� �bm����P-*.�޽�R�X24Ν+����^�d�.^�o��5}����'��Sv���͠��s�6�fI�9��H���$pV[WGQ��<H�@��bێ��y���(J��Cм��&m�|`bH���7�,�w���v	�nЪ;�l���.0i����h}��;�ݷ͛;�6|��F�Ag�SGy�Ç��M[��y���%K鑇����z�ч���*Hx��Et��w���������;�FU��r��!h������lz�G|�|��kojm��*=�m���mQBV|��fL�J�&������23h߁�4s�4Z�j=~Bf|S�d����j�.a�m���"	*J7i���w��e�u��M�."������듕E��������3%Y¾�5��1:���(=�%����̤��8��<�z��8Al��^�(%)Y��L7:��03�F�n<��^�H��ڈ"���=zP*[�(�����34��؋g�!�j�sl���{�f\\ɾR���_�~��?�3�0�&�S}Q�m��Y*�R�a
"f��6'2����W)-�����w�����t��G�K��;�]^`��s��Ϲ�F�{뼛E�,1+��Ү�`�7�f��f����̑���g�����k�Jο���2��쩲JۥSʁ���^ X�`�?��7p�[�����|Ր��%��v�w�-�h� �Y{ݒ���[��{�е����h)�h��B�b�I�1��ްڬzu�h��	A�5Ӯ̖ε��b}F�pgͺ~���SR�阐��(����{1p)mx��H�[��-mV��%�j���uwh���DS5������S����˙�s���E���s,*5�,��x�%�PW��YHCjJx�bY�Plc�զX���ؘۀ�P��WP�7I�̢��4�m�<G�;-�g級!@0Jٍ=��x�*�wn�FT;����=s&h���d�r2a�x�7�ʬ�3)\����4�|:t��X�"�/K�H����21�ʽ�*_9Yߥ�@�3��A@,�Bf�ZԈ�U��0�|�aw�סMg,�Q3Y�����{��`�!_��T�Nl-�B>�Z�uZ��e�cp��4#A��K�_o�mZ��Ru;E���|�Z�}��'K�����5h�l�|�����Y�uO0F?�"�^�Ԧ���b�@���eZ��g>�fj�`m��"*
���~��:�X�A�ۢ˛�:���|=�����`�-� ����O�&O��F���"�yd��qs��\5{zQ�7�@(d�|���V\��a�z
mA5/��NUy�ds���������-ߕ�%5m�����Z�ޱ���>�ڐm�ٔ�]�{�n{�6���fY�	?��b���,<��g|7�!�'�a<���-� ��&'�k�ei�AVO�$V($�)��ً���9�Z�hCt%]᫂Ka�P�H��2�'t���g���ltk[�>L�TfF�J_�]ȧ�tY�0b�ڹk'M�4YJ�Ϙ1��ܸ��N�J۶o�1����]�J�J�o��ƴ�i"�P�v��=��O��[6ӌ�ӥ���i�諭_��q�����R���H����e�;99�

$����C"��r
0P8&**R��bx9)ƺ�gF5y�P,.KymL�)m�3�!�4F�LypMο�����S6E��g�WQRb��>�3�f"�VYQ��_*e@��oh�*���<}�c ��'���Y�����
c��=��ic���8��V�@)+/�+D�-�y6 �VK�.3�~wX
�E����%�ہE�p��5���w�)�#��0�f�y����2�KΝ�:#�������WO��b�y`��F<���1,߳�pC����p ��\�{\zͪn��uP�k��mI�z}��}E��&����n9O�E�E��Z*ȟ�!
����sG�X�DV��-�b&��@4���� �-o۶M�˶o�c�KfT)՚wh���-[�Z��Lܮ��T�%�o'����feA����,��K[g��� O9�$v�ޝ:X�b)hS���c�B"X���[v���m�-B �0� ���
�#�H�~��u�$,�RM�5S^�~���������6�(z��7M�a`œ��q1�A)$T�w����<j�(9��Od�`<��?��(/��ݥ�3l��~p~ٲ��Sz���!�U�ך�'p�SlO�3V�FW�ZM���o:=�n��3b��6#*�bo<����kZ���'�PT��PG�q������j]�c�.�X�)*+ж��?�K��of-*Z����j�PL��Xd沈�S����^L|��꫹�Ys�4so2ˤ�e=�׬7�<p;5z��h��h'@�����jkE�@� cu����V��N͖���_TZ@zk�tC8�뜡z��� ^Fx��$�K�~�e0ϊFOώ4F~[�&|���_(�[�j_I�c8�C���9:��z4r�]4�YSo&C��Rw{�kA��G�A���n�ۗ���1H�i\����}ږI���c�?��}�#�����_�x�������5#�j��̩S��Z�C)
|�A��!/�1��и��
�RL\
%���n��d�==�ϧh[#�Sl|wJ�<��� ��.r66�5��w���'���cG(��7���tAT����$���GQFF�7N�Qa���1J��I�������E,\��F���D��u���O��'�%V~���������R���D�h�ţ���x��/��3��6wX�8��-K�����J��k��M�)�cx	T)A� ��X䥗��ˁ�[�j9w���m��2&@\̱���q0+����\;W
t:A���1lWaT��	r:�r��5�\ap� Wt���b�XC�k�5�fy��_�c�0V�V׆b��D��J�d�>}��3�X۰!�MV	j��v������qV}���SK�T�V<��1f�����b6�U_R��Q��5_�J�@�,�-��鮓�n�M"}���8���ˡZ4,wT�����C�DB�L<��ճʾ�q�|�|"����p	�v�b�<6���;w�D���!�I����� ��w���B[ $\�h7�p���Vy�ar�DY�xQ��0�`|gϞ-��K+7<�#���Cɨ�P��B|�yd��ך5k�  ���, w��q�Fa@8|Ǭ�a�(&f�2�͙3Gf�aH�F�@���^Qƍ�;:]��x� �1[0:1s0�]!��E�d�0��'L� mQ�b�Y�;BAH�9��Y���,<�_��Y�J���H��/���=�iAH �A�'5ز�K�NgY` ��Z�D�gc���5D�l���=�~��|A�*f�Y�֯�����HbP	J.����,�m�GF�,�������� �eC̠�gH�2�����ZD��x���z}��=c�P�9�c ��,�/x����c\S�H�
�,v���#����w��6w%�o����� ��$�0;����r�KS��RGq�!�M���3�x���1�{�x�R����IIt�o�>���SG�o:amQ!�׿��WeH!������?���E��>��s���(����ַ��XRy��OH�$�+�����?�&�U�� ����w"7̐�k���F��L����B ���~�a���~�+������,A��1�mAuFy�p����x�o��>��C�x ��� /�%]Ќ�;"��5 $�{�9)���SO	1���,x饗D0���% ���o��B�[o���*a �+"��F��/ѷi��]��~�;�[��zI���h�P�1�����?��'M��SXF���
�`�Be"P|#��P|��`S 1 �ʕ+� 2ޡ:�= D%L ��.�E�
h��?���3T�b����`�s�d̒%K�hh��{�`0��O>��TpU�7t
A�ҏ>�(M�8Q���dc���W��LE|��B/�щի`���>Vo� �S2E��X�#6�R�.f����m��Av=x�gh���F��E�1���Q\.cƌ�?��ϒ+���p*	��e��U�_y���#����^���>k�,Z�t�����w���� {@�e˖���΀( ��_���?��?�/�]����A �,�,�҉�ʐm �"�]w�%����,��"f�N!FF�Z��6��h��Ǝ��5exI�3,�]mm�����߁��^�_�<� �c��o�2��!��*"� �H�{��7�.x`�+��a�o�Qp�P�^~��H�B�F� �tce!�eC8�/F���rHS�B��@.��OR�j�L�"���{������#�����f����-�V�BhI<��(�q��#K�[n9��%��0ha\��?�fb8A�il�R��_x������c-`A�pb�BK���Ν�=�G;8�f���f��ف� #�����	�.%��f!f��ŋe��Z�6Xd�!��R�l
�R-�|�{��m�AF�A�ۤp��F%�U���j#f�	�D���q�L܋��*��~xq��$�DB�3���֨�����!����V�Q�֣�^��X&5�4f$���7\�ve��Q:p�_@a"� ��q�l�T.������-���R @
b$�Y���"@N��,����ew`O����_�jz'�Y����y�?��j ��7�l��Z��~���к?öE����ȁ���a;�@�X���B��'����R�hФȌ�W(B��q�\�� 3�8��Qf��	�<Ɵ��i�*����B�z�?��ƥ��̺|�S��    IEND�B`�PK   Pn5[�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   Pn5[����N �P /   images/bcd2483e-cc41-4580-b81d-0411c3f5e061.pngTzT�Q���%HI�tIHIJw��tw�tw#�]���J�t�tw��~���e�Y�9�9g���=3��bȈx� YB\X�Y��a����j4�����2<��o�G�Ww ����/�3e%`�QD�Q����E������`fm�`�gk�`co�ṽ�$��]��]\	f�No���-����$P�ɷ)��-%�S1�@�G�(��1.(���4���k�)�,j�����%�߹È��_jcil/�&iBjZL���>G��b�V��q�N;��		4��i�M]���CCC�]���\q*5@EC룕q����M?�� h����cT�����{���H�9~pA�2I�pA��)�te��H�V� �Cvy���������d��7gY�1���{����u���)��BC5���f���(,,�b���F3Z@�$x[��ϟ������w�`�*#����' �	�������~W����P���o�/��ET�Wi_54������=oR�]��v���zMjk�;B������tv	����6�
�bv*(�������}��a��O,�DVL/׭ͶBFC���Wx7/����e�,�tS���`zږ��/1��ꚴʄ��ʪt�-t�4�G�9�ņ<N�~l��VP�[I
�����{�s8���mwR���5�������_�mW���2��v<�S�<�@��'@)r���9]����|��}a�==3��;��C�������W�u���o�1���s�,c���dɷ�.��/�����h���}�OJ�\���D��A��j��q��8S�1u�oe��;������+Ĕײ�����VYul��������c!w�/j� �n���8��n�����1o%�7�n�ƹ�ןT��ҧ���!Ȳ��\���S��[q>�h�rAIY�`�C��ڌ��؋���L���TT���&<���;xYv��A_���Y�:���1e%�_h�˽]e��A���q/wY�/�oE8p��qNf>����֚�%�vhLW��S�����J̫l�%6�_:���FF/3�®w8���]��l<<�W�j�{�fI4+���l���O���J�اN�����qx_%��Cܼ+�r	~�<�݇2����܎GO��%rY������XM���'-,���=�}�vH'f���v�#e�픢Rlc��:*�D֓|�G�!:;��Р��MKE#��L ӄ����
Q���X'�q9ɍ^w��g��	
�l�ԣI���G�5�AW ��>�B=;�
�g��kX�*ƴ���]vȍ��W�b�y��|Tp�JvCG��΅�ay�!٭�hb*����@�d710�޺q��<W�v�><'Jh}G��"�䢃�����;=�:���
=_��(�=�t&8�"�+n*sQ"�C�A�T�t�����U��C��;��?A��h0 ��an36.��w���b���>wc0���D�am=E��`ZR��MMϞ�5��=�`�*	X��j�l�����S¡M���S������@�<�H� ��cFZ5�^@��IH2# �ɡ����� @�������`LR�����t�����p��+4���×����������G�=a�n�����o�w�^�(���'D�k�岿��8�+<'8j���e��	(��opiMx�W�ys�`-D����%��` ��o��y�Oؑ7�Ul�?�'Gc�_5��?NaFԫ-�������s���I��ߡ����ݮ���a!�	�q���ߖPnl����G��.LL��7 cɫi�!tu�������J{ �F����WK���Mmږ�#�ص�TE��ǵ
;��2Eo^Is;]k�'��Z~���o�hg���� a̼Q����9�a���,��� Ɗ0r������g��X�#�#1�v&�U���V��/$d{Ͳz��ܨwEHVF�p���ۿ����9�rKW���WQ�D��k[�+�W�T^��H�q" >h�)�>,j�ZN��ߐ&��Jhn�.ZB:ނ����Zvi!�dz�)�"�J��V
��Wɱ�:/�,!�՟mO�)��V�ε������D�r�P�x�	)�1����kϤ�yhvv�󗮗\�o	W	] �t�W����o�0�";{�ۙ��[��#��1f��W%���!a&ƅ>�U��h��>��&@�����*�+X��[�f�jq�?��0�_��-���Y39Z���c��ҫǕ��$��=83��P���7��`-��
ZY����J�e��t�x���.��}��#V��9H��-�gB��/�T�gl�Q�<��� ���M���:��T ���A]�fYԗ|�K�k��� �����1���x\4n0+
<�$PLe���E�,*b:O5�W�d���<�n������К:��k6l��'5������a��]���t54�^SF��g����0zv5h���M97����D���"́�����Y� �[�A��a@u��F�s�θq܌q}~>��?�6���C(����,�TԠ�Ł>UG	?�4�������V��/�-^�]@H�?A�����h`��}S�Z`!zx���B�r`-�,\����<(�.A�#T�5o�_c��k�B�O�) ������������� s��ScE#A�O�J��Ą7�l��{S�'+ȫ��<�\hm���|�2��[�{��5����O�bW�����ў��@��w\A���� |���Ҁ�T�#����4yA[���j�E�����:��ը!��5e��cy�`��蝹[u�yN�n�4┬>�X���!�
_t��-��aa:�nF_b_n̶i02"��ҁ��B+������ρ�F�
���dqGډ�hl;�[-g�%��e��O��@��P~(�Ї�ĠN�ɜ@GO�"(�[H�;H[��uܛ.�O�c�oeu����b�>!+!XKS6~L�ۯ�1eM�h=0|whOl8�j�`�ÈZ����^�)�6�5���_�c�*���#���u�/Zǽ"�^�p���.���L�ľTU��������d��5�1Z=����Y��2[����G����͠@���$i�V׏0 �����\����GT٬��|<y�Y#���C�aG�7X��fiO��Cw)�κFb�$�Y�IB���2iM�����Q-I<��.�S���� ��f���T��}��d����vņd�~�<�[�X�g�[%0mمZ7.]���>�>LS���Vn-���םh,so�(7$%�a؃���)e��1��o�â�`�ٞ.�YbJ �DN��z�J0��qGY���m��:�n-39��P!U`��)��z��y%g8R���<�����40��#����yr��O7�$�(2�v���/�o�;���POxDP���{]k�v����#X�B��T ��p$Q�y-��I�Űr���>D٠�"����,�3��>E�x�!C�@��E�� �8�k�r�Y��T�|~�c�{b'sg2�eG�"K�f����1��fr��x`��������a�kSs��M$.�]6��1#�c����L��]�o����eq2��v��1��z��!�?�<{�R<��?�`��$;�c���;oq�#A�A���!��*LE �̬�/i@��˙����ɻ�B����*��P��=3Y{�A�R�k�3GF���zPM���謁V�N��/谵q��2��O�G��'Ԋ-b뙗�%�)?�ǆt���1���Ȃ�u�m��C�f�KL���k��0Б�&���G� 7�`��+�f�̡�F��WT�y�t�l�A��||�J��i��L;e'{��9�����͝�fG�]4v�%�O���6#N��:��S��[c
=�uM�\�+���%��[_ȟ����-���Ȍ�t*�Γ��Tn�x�p���bR�K� w�w[�'G=�ٶ�$Op � 9�6��F�#0��6{�����Yn�J���E��1I3���{~�C��>�Y���r�8A���]�D�޳�1�=��&�W����VAv����'�#	�2��h��|l�<S�%K*�
u�0f��Rr�
���&��+��"ĺ
P tl��_�5D�eTʉ_�1�{5!��@E%���(�	�D�s+`�ǉ�E.�nU�l��R
i+%E�{�2�O�(��\S�&��,�ȱ�%V�>1�ޒ9:�ѮV�}�Ҟ��ȷYԚ�X��+�!)QokDX���X[��\���ݬ�أ��V]��-�1˼>�Q$�#�ñ�@r	� ~CTd�Kl���2��SK�A�CٞV��.���1�ܞS��,�Us��J�/�^����� LR�^��r�`�F��F��dK'R8�sWdE�#�'ȋi~D]��hd{��%#�����^3w�$Ǌ��O>-Ö�3ԏM**1<�2Tc�m��P��;Y������v
�2ō:ӽ�}�Oq"U�?���F��U�`��X>~o�R�E�1���e����	]���<����+��aYAU	�Q�F�?�@�^b������,wMb���RCY�#%�*A9�Y��Kr$���0�YȎ+ ���ܷ�VO�2��aw��2��9��P�8�g��-�КΎ	&9y<H@7���R�/�/i3(�C��ڹ�/�N�%��1�:��i�î�����$��^��?T;���Oa�C��H9P�̰�eu�Y�Q5��2j���hl)��Cau�b��o�~�Qs�@�%����^�����bfJ��~HI^N���+C�st"�����]�l;�"�ث�s�n��?}���E���IRY wG�Y���Cb�=!#ຆ.�FR��јf4���b�2����Ao��1�p9����m3Rm�v�����2J��q^3>BO��}+�X�z�vtʐ�7��ډ&V������4���k����ؿ��E9�5��q�%[��J\��T�+A2��q����P`����^����C����70���W�� >��9�9��6f8�&m)�G���%C����Gf����s�$-(�o���=���cJ��,hp�
~�����zS�~ysX�@�Fū4���t&��u�0��]��Iu/�xA�%Q�j�Fd6i�/��<�gL�	@��RD^b��B��S�&�TP�"�c��Q�"O�&N?���
��)Iy��7�(�%i"f�][�؋�ѝ�=h�o��}����,Ӌ��&���T�r;���$�����M����bA���j���{�	�M�_~�D�������NJ�%����0:���� 5�f/%�3�,x���]���]�d�G��{��P���c�wP�gQ�g�����)�7TCr���\���c�@�ʹ�,W䴑�n���=��g�*��t,F�5����rL��T� �i&d!�+�0&t��+�;2ߔ��Oò��'����H�
I�y1��#K7&�n�)����F��;�8��-u�m�b�-j��&�ȑ�Q]z[Nt���[�Z������I�Kޭ.��HL��쟔���
���W'�6��10Nt�PsM������^n}�˥|�vW���۲��ɵ��7Z6�1��a)"0���"�l�p�Q�2����6N0���3�����ֱ��	��p}�q=1�O_͑����08�R}�
p�9�"��Z{z��U�NH�]���~����'����{����Mb8;^O�Y��'�0B+q��CJ�Ž#�6�yl�;*j|{ɳ:	 �b2�"}�Jt��@p����D�ʅ���e4UO��2��o�wX�(P���������2n�v�\������K�#{u���un�H�Y���e���ؠ����l�%�}���/��U�2�{�0ؚL�����^m�M��������!GѵL@=�Z��]�&u�I�wK�"��fj�hU��4d��Q3/�]�A�h6ȷ��|���OA��oit���uxq��� ���kQFhIeH�ꉿ�DbR���L�P���VP���ѣɰ��|����dd��7]���Y���a�0�57�ؗ��v5�$��Y�Ϳ�<	mQ�y�Q��N�tI*&;b篏�%��)�)�Wy .�14��&�@s-N2��ړ�y��΁ 6 �������#��TĀ��̛�?aG�V����sϵ�l�)��b0���O�8��{���u�ːp����,CW?u �2��Qhf����ͼ��PI��i#���k�T Ѐ*��x�,B�ϐ/��D=ܻ9�_D��	�h�]�O�D�
�;�=�c���Nʮ���;��'�����1��H�M��I����(}��0%�c�+k����(�_�r�ɧ�}��Rvi��&=	��W�R�~�DD��Za5�����gȽf���������9?�O��?�8�q��=�%�6V_f�$o�=:�ÏD�|�
�=@Dz;�&Z�n�h]�a����v�� j�,0ש��o���
a(]������B'�BO��R���l��j��p�-�Rf����=D�R5���:�1J2;	� ����/�FzZA_T�yO�Č�\��TT���뽰��TFؔϷ�B�nȫ��K�"@1J��Y �dis90D�y��?�Bϑ�D�;o�K��~���V&�0�&[Zs�G��.�u)����^�0�t��xj�+!�;�h�`[�?Ԑ���1<�O��E���`�t*��~"<��y�q�Z��K�52v�:3_k6ab�:�T��AպD��?�V�S�����H�U�G��c4̩x��'�}qy��ڏz��T4ڴ�@�����"�~��)�A��]���b�1�lM�Y�ˏ~pxW�=PeE�����n�]��5�b�w��fT�M��jd�&���!-$���R��{�N┕;< 9���H�	8�
᏾ϗ����n��,9�p�����"��V�����L[p��@2��̐P�Z��ΰ�8J���p�����.�!U��"<��������;����	��ܛ�/4�^ޥ�Xv�JE|cl��`L~�Ӂ���|�"�KI��9��i)}����vl�)����5�,>8�3���=�q6��;��U���W�(Cr�\��ϹyR����qx:5���|�Zw�VuÐ�s�J��$��/���5hxX��8"U�xF��W=�JJ�;H��JpVm��}"2"E�~$��'i�/���ܴ���P�V�E��C���zN�As�=�&��esK���l�lW��f��hM`���s��ޑTn�$���2#Q�|l�z�d�����)�ȡ9{�&��cE���"���o*$�܋�n ���5I�f-��ۺ��g*�B����r��-[6�7�'�_jOy`����R�M3^� Χ�l��X6�H�����z���<�}�EG3 c�Q��<u���R� �i��م�m����h�����b9ًl`��K�h����6�Ɠ�Y��3ךJ�횕�ԗX@��u�|WZ1�;� ��v�������k����p3}�K�䵋������'Q&`�F����%� ���V[zZ���ɧ"�?C2;=_��l9���آ�i���)�6���R�h',���m1�ظz����/�g���WZ��Q��[ _bH�7τ�L��Bt����<��G�iY~|�l�����d,:37K��?���ڍ�-v�t�+?�ȼwe����6��,�!h��������K<�Z�P{6y���Č�C��~Y9�'���~������!)��m�3Wu��b2�V���%߼k���AVs�K����꟔��^����������ĸ^N+�%3����I!<�<ʙ�c�תA9�����<,'�ʴY���&P�[3x����|�VW1z��U�H�b 9Zq���F��d���rl�'���ǚK���JT��1Gi|w���v��;Q���KŮ�b;�ҭ����,գ)s��_o7�.y�5Tt:��˘9�_;�<]�ܴ� /.��x�:�W�dǡ�JJԿ��~�M�F��JKe��W{�z3���j��氳�<�as��l��V���fg\ '�9���O�7�k��t&<2p�W���x�/hvm�I`d,�Db����R.����8��bjr]!v�g?��6��#����Rtȝ�Lq���jd0U/a�z����dm�	qsg�2��J�ic�C�o���f�ꢟv��0�-�ȏ�i�˽�|td�cOA�o_��p2��4Պ��`��4��aM��:#mD�6$}_���{6�Y�<�@|cY��Ҵ+�f~P��	��|�^2�tWPh���r���@�>8b��
a`.�n��@��D=��&b^(9;�����YO�����D��92i�h��z�e��<yd#ʑX����.���wy/��=Ǟ`{��ݱ��I�
��?~��f��0�G����o�^�ý�����f饃��i�xԉ �Y+XT��K��6�/��e��V�{ً�x��H:�(Ʋrm�rZf�����+�n55��I���.�nf�ooNz��D�޾>ׯ�"8�oLl1>}HM΀y��X���}��B���S�5����ȭ�O��Ψ6a+Jz3���zw�.9����������ڒ�Ĺ,�P�uZ����B��ڪ��-M_cT&>Eʵ��-��%�ލ�
]��".D���5L�&m���V=�Ӧ�x��A�0=��������x����jgC���	S����N˹�� l6�"Ƌ/�������.��K��=`�0�A�?�D;� 3��P6���,-�黡�,�����$��5��l��O�-��-)��{l�oJ����4ꃘ�Jpm竏S�#����;���l]e���1��BZ#�B-�c���+ר0�wwx�s�g��&��Wߛ�t�R��=��t���ȧ�=�V=7f�&�d�a�y�Rc."+�w+�t���_\v`��g���d�sg��ݡt���"�t�|8Y�y#�/?�$�i��Ģ�羉�lH���^��8y9E�S�M�A�f��S�O�<B
��n���?�6Gd��àH
E�{%�?&$�X˘����ǧG$�r5�ق��:hR{K���O�6��7et��㶢����&�ک���e_f�Q��ގx(HJ?m`'�OW�i��a�h˃b�A�\a�g_nu�|���]��|� I���R����H���ʋ�mDY������4;�c����5|����f�e�s`��q��w)�lj|��~  Ԩc��#�Sz2f��O�"�ř�9�����{+S�y�@���9֢A&��C }1Y����*����4��l �bW��#�sL�`��N8Fȿ�;��D�Fk��2Z�I q��w/Gl<����6q�Le�`�3�k���������5���o�>��oS��T�ֹ��Vq;�5�$0m�+R�b;3<]��m�+��m�u�":�;�J=j�����C
9����Z��p�e��r���?Z��E��Y�3�$�a�K�F�e;�U$;;�;fxLQqQ����B��/��a�s�)���+�e�W ��B�:�ނ���f\0�qZ�("�0�s^j$���U���ֹU���Z0���C��%|��q}0;�ˆt�HS�W�lʀ!L��-�av�� NW�	�w�q�Z�����Q�I��˘U4�� I��-6o�s5BNX�b�6�8�4H[Wuq/y<�fT=���}���{�D}t_^�}i�Yhg-��X�K.�4���:�Q
.�|�A$AU.���#���P� mۨr.Ң��h�GJ��+���1x�%�:�����7����5ג��8~p� ���!�4
MI{�r��1�:>eE�,X���?��iT�a+���v�BZ�?)>����df�mR6��O����ĻU�#KR��6��-s�V�@gY��c|�ձ�I�6$��Q�
�H^������gio-c?)����!f;K��}C]p�۔v;���ϟ��p�5=\~��X��۴h���!lԧ�?W��/!�Y6��6��Wⰹ=P�&�E�E{�V�q���4�in�O�w�@���mC��b� �Ȱ��<d��H�~u��D����=^s�/avg�!�<pqOLÔ� �1!�]U�*5� �Vf	��l#:n�NS�/ϻpG��W�k�T)#���Dv��J�`3��WĽ��>�W���� '%��Yg�M�_Ǵ}�B��&ӯv������\�nJ��y"s��&g�+#�0�fA (����߹ߐ��EeQ6�Z�A3x��%��V�ܙ�&�ڙww���'j��4� ��G�a����k ���fXR�I��9<�Yrn��R꜓�ӕ���f�$-��6��v�6�h�G�ȃl�5
&3���!Z���~Z�tF�ν�bm_!{�Po Y崅�}�z�T	L�/�h[3Y¦
p9Կ�q����Tjg�;��T�,�EU���%5MB��~�mb{JJ������1�d��[� ��Z�c-���(`�X����hc�.������N��ޘʖ��ȫ�R[�K!�������B��Ϯ��/����vFU:��M`�(�`Q��� Q`��T�Ŏ(_ �0.�Z�L�R�q�N�e���ۀ��,�X;�,5�m:��RCT����ϵ�k/��)e�.1+pH����ל^�l����!<�D����x\���y��OkAi?K6�*39�����W�A���T�˭��HZO7�E5��|�Ͷb�Ef,I�7��i��W�. ��hٵ̥䎢�%�;I?w�~��ǩ���	w��o@��$�a=�������q`gf��|v��-Bd����v[�A�2��7Ā��g]�a�����T��qK�@��������v�����W�A�9����(8�2�=�	�a�
��+����*087�p��c�u�Ⱦ�@2O��Nqe"w�ǩ����|l��
R �'����|"i��
�(�MPA�\;��}b���r�f�]T^��F�d4�'Ŕm�3��q�H�Q�*3�H8��އJ�C�\-M�n��@뜡HHAy�#���\A��$���n��%H������-t�Yc�}Xi�(}<@}���pfÎ~uI&yk�@�1����Ј0f!����$���[����.�6�ACC�W�llP.N̖�Z��hk~��HHt�
8�SD�.����#R�����$�a�DT��G�x<?^�8v*��M�0U,(jv�l��=z0��X(BQ�����2 84��5W��{k���
=�Ͽ0l�� ���PM�_%������5���=����a��7�A�&�a4,q��&���UJ�*qSjT j�o]�(�y7#��x��N����M�#1}�U$�EH�����(��"�X�92ι����]��ɮ֮)��_E3��dWlr-`�:��%�:����E��\���!J��>^��m���:p�l4���� �;��q���C� �8v��|$�Ϫ��ˣ����:	��=A�+�+3-'^��ơ$�.ى�Q̿�@m�DM�
e��������P�x��܃�Y��������F	Ҟ�X;�������ƪ�=��Y��	��o�R�{s�-#P�|8���"롆F��	~����w���ao'�^w�c&�G�M��_�#��u n�n8 <���34-������;` �O��{�>�8Jߍl/�w1ϰ����U���p�!�_�3�smJ�{��@�+�.��҇�2�fb%0W�#V[>�28�&�|X�~zíI���͉��n�0*�/����9U"\�<���蚿zz60ے��S&Њ�������O����P��Qa�=`x��@H���m[�-�;��os٤ͭ�ΓZ��=�]p�k���Ny�v���4$�r��r�RE�an!�٥��n�k9�Ѕ�iMr7ų�3�.��/\�n�%���9؈M� �����vK98Z���(=3��� �)�
��?�/������՞��{j�ɸ䗋�>�O���f�O����(��˼w�6Af��_�g���A���j��ł.
�Z����IN�	o��z��t$�2�����e��@���Da�MP�<�󹂌$HN�3~�HD�}�E!9��YO��Ǹ�fg��]��YF,؀������R^3]������Ӵ��|ǋ�r�\��sf����M��=/��}��<��nS�~q���To[��{}C��R>"��\��I�q+����i���9*�LĹ������*4���LǤ�Z$��֜{�'�ʟ���;̮���W��̟����źK��P,:l�}i�9ig.���(��(���+��h'3��gCl�i:������6�f,��d.h/8B9θo���c�9�Ϯ$��� ��ER�8=!4_63����� �+Y}C3�Qh�^�Ϛ���沫'X�5���O?�9�N�� ��|'KE*���>�+��G_�Pcr��s>�8x2�n=O�ip�g��"gӿ9�&,�N11i�-BʻM�)F��e�$s�A��4�,������>����c��|͖/��|Y0��Y��M/k��3UR����ݰ�lA�K�������
�vd��\��[$�c��R.9r������F��.ϗwR���D�_�~�=mu;�;����]��.���-/"Ã!���s�>Nb0��j��EC�p���(�l����d��2]=<��Q�?�I�|հ���QxQ���ׂ�yq�5rBY��������B�Ӓ�g �%i���1�����cPsf�3����p?߶��]���@�H$D�ZSr����K�
C��"��
�E\r�?���]|Q�7��sw�9��8����`8u:p�my5�1��q�|5­���fi�@v��G���GT�v��]ˢ�@&@���OH�	�B�aN�d��V�WY�����.�����@�(H�+���o����G +���zϚ#Y�='>��1a:���kz>X\�u��x�`1��\<�����M���ơ
.Q�H)��0/��yѸ����/�kq�2x��XZ��{賏��b���I%F�X���H���{#8��jr��טK�?A��U��/3�:��Ly��}>��u(Q�M��!�/�W;�4���]�!�H%�T�%��}o;"�"��[
��1�gO��/���|Ԝ�}PP!=c)
��ߓ��.];zV����ǀ�*��d�.�ϕNM{~�z-,k>�l�%���L�Y�2�a���-5,kF�P�H����~©���k�(��Zyԭg1}0A�CS;�]]d����L{���A��x��#U��%է�P�qS�]]i�����+?���q� ���y��,����W�Z���u�-c	�N������\� �]�>]�|M�PC�N���vWl����Ez8�w�Pқ�v��d��]t��	�\1�}�I�������:4�����P�}EΥ԰�%����[��j��D�)ٴ[7�a�z#��uB��㺲H�>N�8 �,;۪i�>7���5��gn�^{P�RՒ�C��ڵ��d#J��s^Ђ�J�s��G��q!���O�ZURN������.�F؛�Z�v�*�G�o~Tؘ{uF�9�LM��,T��}�E��bX/����H��0�2�UWkmx���d}2�&��)j���Jc� z�iR-���۽_��n*~��*4���t1�jq�Xꋣ1��>����oA]Šؠ!��"|O�Z��1 �w���Qs���9-s��.o~ƪ� {����w� ��"���!����٦�i�!���+mWKk��6g����Hz?W�
[��c ���	,%Ѐ��&��,��gRwJ�5u5�8�&5������a�5�f,$G}3�S��D�X�gU����b���೘�/�w*��1�X��z����<2B��?6��?�=/$���s�.j!Ċ%A/�\R��x_�|=ޑ���.mJ�`ܦ�f���5W�)�l���GajLM�5�ҋ���Ma��}�B�ߴB��Dl���g� !k�+�f���{��=���S1A�^�X��Z�]V$��]�Ar�W�I&m?��א>��j�^J��B��m�<���C��-7�x�y�%@�����9�T[@-��
�)U'����}�u�8��\�i&�J3J� ��m�(x��<��ySKX�7!�>�|��Cp�J1[��=�>��-JE�e������[��f��}R&�n����GNs��[���7%�E�5��K¿����C�R������]?ҏ�����h\p���������˲� yr8����6u�/M>���xe�^�N	��s�OW�#.��>��]����t�M��2D�#�^+���1�J�uw&�yP�y#i�l���t�LM?)Ws�X�v�7'�?S펫�9�/j.�6�U��=�"� ��H����pӇ�ȥOq�w������_Z+��L6�hj��g�t��0B+=F�'t�@�E����<�5�mwMޱZ�z�����T͠ pL²`�� RCL��S�b�ʁ�e���./�?�f�R�d��������6R��&�%q\(�f���=Q��H�;�O;��`����!��Z�~g��� x���̮5vg�=1;�����D�
��'z�	����*�gHI_��?���]n�8������{=�����Rp���-^j*�`t7�����D�A�w�	��[�)����y��?����q���'���s"ɋ�S�-�W#���@�O+$}?��o���)��j�[��cD0�,�F0���D��(�q�g��;C��'�(�Yz4�V��z�q���q�>�޽�{γ�M�EkNͮ��7�(��Nj�WE���O���3�/���@�|�'jF����K5,_j�Q�ko�>�N�5�R����m7��}�,�Q�*���m�2�;3�FE��fc����^<��9�])Ex�{��7o��I4C��-J���r��D�)ƴ�e��4����Ei����i.���N	�G�É��z/�9��z�����%w6Чn��Xv�r~�!�#�9�M|1˭�hp�>�i�a,FA���|?�}��އX&Q��š��տ�S���9� �^�?҉���8ʄ�ߛ��	��Ԑ�Ǣ�Zw�ē�Y����Q�!xԀ�P�o�=���(r�+ ����#
\�k�U��L���s���,�*$9[iFYU!.�A*0�( 
��3�9ju��+佃L������&����'�+�9��JЭ��z�Ԗ�i!�WVN��?^��+[+�y�32����q�"��(�t|���F�E(Ñ�A����4��� ������
�BA��/~O��6P;@,�ΨN�c�쳯�~aU�� �kr���������!��m%l��Sb��F��ŴJz��Ҫ����}�6�2��Y���F�2��c:b"�*��6F�G���3�㱷�JVA�jN�0�����.K\�� �j��6���o(9�g�~�|�5X���'Ca�<QVC��X��l��j��@���W� �,"f��«:��4��+=�|����)��zF�+���p��Ҋ�=��NI����Ǥ<���.�Jd�ȑ߻׬2�F~�+zP��W�cyOɗT�y�~�/3V��O����J����&������Z��`�yv{�]�%���;�R�� z� ��j�Q���
>������c����}bQE ig!�+A��"V�"��DEFs�~�Љa. W�PMjN��]&�hVr�'���@펝�~+�u\��e���d������a�$}F�c���p����H�V��d�Y�\�i��]�ȴ�COBY ð�؏�t?��C��> �gU1�'���Q*���އ@)È$u�z��G�Ӎ&��ɈOBg����%�b�C~P���֠B!k��G�VL��&,Ԫ�E&9ٚ��)�0���l�!��#^l�����N�1K�9Z���(��8PAkj{���ԁN�ۚ�5�A�hp�RQ6wŏ���W��w�4�;͉UZ��g6B�]�v6�z�G:��lx�1�$��Ҟ�0�gm�-r*��	!�d��(�V2[5�AgZ��?���:{o�q�]�h&���Tb�%o?��`�/f�Yf�O>�g���8O6`�O��zNn��$�? w� Z��d�X�O�dt�����b�����  q��2�_�!_
��IƵ�V�M�[�viY��3��Z!G{��}�$����.�F� ���5}��0����i/��/�<��;U��)��#�4G�aCNKH�+�0��bmTvc�i�|��j�'�����hl�ZN�}A?Y�o���X��z���ڳ��p���d ����k���\㥃.[Q�}$��G}����	o�-,�鈽s��vu��/w��/8��F�(�tϿ�+u��@����x�� YHT��UsX!K��'�v�I��� �
04u�y�)U��|��LِΔv4�X�`���޽�BF��*��Ǻ�O�F���--#r����e>�O��vYm���qB�-�XzD�)f�p�1茧t+�Z'6��Ζ��QN�pk+OG1�.s�1Sn�\h��^����!�0��ϋ��.��X�Ǖr��\i&vN9�\:���{����UyPq2��-��g��yDm�nT<GN��8<�$S�8�h++|�8#���8}	\zyj��8��C��M����뙌���O�V���v<�w�\Q]qľ��{�rf]=�v@	-	$�����Fr'B�C��+�����$�5-Ѭr �ki���ԙO�z�܆%f��y�s�z�}�ɺ��$�q��|Aa�i�:JG����d.ǒp��EСr���IB�'##Y)��a�v�!�"�E�"�?��: �7�.!�H	+]�-�%-ݱ�t���4��4"�t�t7(Hw������{�ߝ���ƹ�;3�n!up����.w<�o�������x {�@8M]ӽЉ/���u��g{����?:�Q��g�5��?*|�F)Ab��N�"�N���PHt�y(��?��(�W�XS�{���+�@���)���\�F��g��q��z���w�3i	xq����]���t�>����Lk�@��:F�t��?uD�}p�[(��U��#it5�*A%�job�d�j��c5.�6�:��=�]Y���s��hj��i����*��"<���x�2���&D᠇�_�S׋k�Y���D.��8@%@����|ѕ/�+�*�3�+��]Ș;aRc���xP���P���h�3ϻ���L�YO���ׄ��y�B���3��~�8�&�G�
7���8 ��I��<��� �9���X�M4��5k{RA�*���e3�O�\�UA;��$T�l���V��\<F���i��ţ-���Ww,ZS9wbÉ����F��� U� �����2&��'��ݓc<mw��D���,��+�m�5ma�f��=m���j�f0��lԢe`ȳD�����V296$Ac>���Q?�{n�X%�r���0�>N��G����zO�vM�#z�D=�b��� ��e<��:�z���а@ �-Wu��d	��@@��|���3y�?t}�W�yj`���m���Q� ��'�U��s y�o�.�槮��)��,�eQo�ad���ڍ
�]�S�OM02�P;xM8.��':����e���n���3`�*�L'q:��3�	$��1^1խr���}/��&Ҩ �L��B�k97����y�B+�y�#t:��K0��jNH� ���)gMR�lN���p�qt�m���`k�-���?�y�`��B%�-8�ՄG��M�f&m�O�%��W�<�����$�Ze��tw�x��F��| � =���䳡Ɛq(k�#.&��]�J6�*!����0�Zm1V�n+��E�t��� um���F��j��l� ����XU/sV)4��k���x��;�$���_}*���=�����f���"��|�4�c�/�.Y�X'<6q��n6�8�$r������t�Zqf$O#ny�߷@!41$�,�~1E��$B� 3-q2����I�b�Y(��&ccW9w��j��a����u�����a��*�ҙf_S-�a�gaذG�wԼ-VZg>(��{B�1��D�.�L�Y�KV�Ι#��t1�������,!�)av�!���m�U�)���>�-�Td��<�xJ�uW��]1��e�9> �M�����E�y@1�P-�KJoeA�@�fM�Z3��g4Y�,䱠 �P��g�d��&+F9�����Lω�K����j*�l�
�%C)�A-���jx��X �����egV�q��КG�!thl|$z�X0e�aSc��2݃�t'N"�H\�N��W�� �(�;����Xe]������Ն�(���0���[�]&BM�A5E�o9?�Gtlz�_��Q�Vx�,�95!;��T�/���G0����t���ƭtOl<�`�pػq�����	>JdԊ�w������,m�C\$���R��`z�?�C��M0�����B��57����?ۙjG�40vz�)w$��3e�/�A��
6�x����)Ť�TS1U�������������Z��@���X6{�n	��4��G�S��YJ ��y��@BtG�ۑ;���[��u7����NFf�ȃ��� ��Lj�޹�ˌ��-F��R�7Ke�տ��C�������jp�ËW���Zi����>�)u-�T~��.��<t�'�h�8	"�ieR�vie���oܥB�j�w�J�f��x�$% ,�󵥞�M����w�ߝƀ
�(j�m.���i��@�j#��x��Ž`v���S}�a?g� դ��5����F��Z��q��(:��C��u���ڋs�.#�3��H�Z[�P�a����$'.�k��ęB��S��i���%��������3)
Xd��3�P��R},�e��8������Hu%����nꢓ0�OZ6Ҩ��O1r���/B���W�ٶ�����$���s�52)IP+�%�� ��G��r���k��*i�{�����>u~��Uq�X]�۪�EP�I�%�1�WpI;�4�?ha���R-*C$��ȷI�[�mŤXډ>��v78T��җ_�W��`�ǻV�o�~�%�|?��X������	����&��Rn*+KF|a[c/�g�m\<�����2Fᄁ�ǘf���k��0K�|�x���ku��5;�<q��A/���D� ��ԏ��0�!��Ж��U��g�mc`"�%��伪l�1��pT���w����I`ٿ�%��|Q���B��\'�vv�j)��)�;�#~]}�W=[��ms���%PX�W�y�{3'���&���� ���f�G-�?G��(w]��������Kc���alx5�M�#����H�'���*H���w	0%��;s��y2�l�$a��Ԍ���PB�$��<�	wm�â^��X�k��!�vA>�� P��?Ip���PX\b^�){��G*���x,>�A#v�-�/��	���g�h�-��i�pG`"�c�����R0b�}!�l�$�;�+X��Bu�"/L�fB���Q	#�i:�%�%Mh�h"�"���u�4{��[����W�ҿ �Vd�i[���0Vs�H_��γ�%ח�>m�Z�=�ͬ2��y'm�����3ۡ;0|�p�������׉���[⎤��p�YJ���:��ꜝjZ�ߟ@���� r"#�Q��~����z�o��g����w��v���V�I����E��˸5O����ڝ���M>m�N�g���0�h,X���O�ۢ�&��=IE'T( ɹ�b, ;�,��V��A#l@�j�Z9J�_|��a�:?:���*t��"2�C[8���=j Ay@Ċ�6JL@�#�QfÁb���Gy�ZL�p�9;�!�$���}�HX�Iv�T��x���?����[ k|?�c����b⬾C�������Q.&N]rd~�J��*~dA^�5�v��J���4�2A�]�$������
�F�>�Er�IG��Q�S5�}W����XҜI�˂0K��x���Y*L�&v�x<�@�Yu,N�ہrA��)�B	�v���᯾]�Yt(feF&#��"�<�8���tJ���T!:%��#��ҽ�n��Y�a!���E���:ȏ��o�����{�Z�Re(�삠�:�L`�`��%����\�|��:/&ܟ'oƙj��h�ԝj�$�fJ"k���z��:�_���w1�ш}4Z<}Y9f�5=e最����3��uWG�\4�}���4�;|�����Q�_q6H⠣�����.�p/pPt�0�尠7%����F��Kn���f��?�	`6&�������c�Xf}*�D����μ���R/}�:��ޢ �QBջY�Hj})?�h��|��|�ł-�AeQ7%.ep"����Vxx�(=�;��~y\�+�/�@���_I���θ�[󯲚L�-WH�ݿh<�B�7SP�z���-̿\����<�2�0��52�?�ΤL�5�^!q�P�+'��U�2�m��r�o�hA�H@J��-�MG�sV�ܬ�����Hi1�iX�H騒�0�u��O����i�)\�L�Oς���`�kon&-w��_�k&WS��E�����f=�U�A��0��)nv{���3����n;X�L��0B���#(�^g�� 'T֏ ���a���6�hz��g�+�|Y�<N��q���[r�F�R��dAM ��L�[8�1��?�p�%c&�+ɿƕ�,x����>�x���c�:!5l5N���^Fw��̝&��A�$�,�MvwC����d�Y<gaA*���`��W���ّ2
G�8jL����ظ=�eݟh��2�,9���u���w�K��g	��8�M�J̚{"��p�ۗ&	�?r��0��>S ���uq̄t�wR���Sm�s�`QVnq��h�Z����5�Z&�$����׿�.�F���<�gt�}E}����a�ς��\��	v{�M�+���qgY{����3�鸃��g��]��J�ӁW��ϟ��ښ/sj�N��փ5���S/�8U��TP���Z�J�Z���(�NT�����C���J h��~��FH[N�}8�PtR�B��C0[����I��L֬������!L�=�hI����M�TARb��z|�7#����h�̢O���I�_�aX"գy2�G~�j��b���1.|n��x�k�wz֟�$�J9�	Q���]'���{r�?��� ��?B���pT3M��� 0&�=�y�S�!�՟��0�f�Qq���B%��(18���k�!�sE-f�v�{��q������HZ1��Ӊ� �"l�!c �?�,̵TK�D_/��B_�rf����8]E[���E�ܧa�r+z9�|�@F]I�z
��9( ^�ŭ�[�C�o�XH�t����7i�$�(��V�b�/z�i�t�����7����vi߰ێU���A��,x��Ր_�H2��>Rӊ��q�(<�*�� �!�&2�6P^��6���/]��KA9�x�4�t.҂�= �o:��za����A�ne��G/@k������N����0Ι��t�G��������3�%�_�B�TTgB�sj�^ �I�S\1ѱ�Ӌ�`�u����A��۔$~@���8��q���{^R�cq'�� ��Jx�&t�. �u�Fٱly��ɽ	Vn�O�@+���������ף���5߿D	�%� �r� NJQA��#t�n��K��0��H�E�y�VQ4 ����'i�F<@ɤ�+�e!�*H*Y�^��&Y�����0�����B)���9A���JV��<j�R#6�[��g�J�}7�����)M�{��^Z��v���X�����`�%��x�n�����+{��Z��rU�[��9�<�9 �W��(� ��� ����DewC�2��e5e�	�XR"���G��{\Zw;�m��4�!�^��� �W:C~�5e��I�EJ�c���r�B�4�o^T}F�� ��t�9U��=�#ta�z%jp`S\@LF��O/�w��9(5�d��ϫx�Pm,�#T���{�c��Ko�y�쁈 "���Qo���(`�8{~�������������_�0%:6-
����v���	Hp>,тwJ��Q8�V��*N<>��I�g-�QM��*0����8e�����쳳|�>tcB��e�t�1&�rjM���3Y�pYB�8~�V�ϊw憇���,�^���	�#Ԇ�gc~�͝�9�͈���U�L���-�I�a[�
0��v�X\�,1&GTSr��%���B慶 ��|�4��E�ɂ���Aq�8Z`J��ђ�Zc�uLL�[D�"@hT�I���X��~��ڹhT;����jEw9�Ek���f�e1&��z���D|(�Sb�УR�j���ڷ��8���>���9*���S�y���w�����T�Q�̸z;|@�t<^*�#�B��k?Q�Q�Ce^^kEΛ�_~�j����U�����Ig�.����s�͜�+ KG�̡?Eo�7+�=�ei�w��越R�$�@�T>��yR�3#��R����+P���x�!+1���sz����)Y� Ӑ�N��B/�~+	��
	h<�ɓ�����JMq�x1@S�3�I뾶�}�w���+p�c>]�ST�p�3 �>�ږԦ��u��m����L�2XZ�ΐ�Y	�ؠڌ%.�D�o"c���x&L��e��@�>���������O����\3��`��Y�N�����o�������X����=����$�b �̖��nX���?�@2�	�=�@RM`�"�:���[�؃eSFw_�+�B):�6_]Bb�-�K�F!��3\��C�D�F��֥���/ӺPʗV�l�q��σRS����'�1��qy2�V8e�'�.���|bbi|���;�pbF)��}���=̀!G�
$����p�1� ���x��逝4��Z�p�v���V��OE�$!��l1�"������`�?Cz�L}�^ā
⭱���AΙ�I�D:�m!�-#qF�a=��̷}[
�I�� �K�8�T��{� ����"ژT�<�Ol�b�Uq�p"��Rª�.����1eOfZ��N�HƄÙ�Uڑ����EU�D�T�Z�Z1���f�T{���7��]�����-(U���b������+q���X�lq@EK,�P�4����#��,�ءC�9�#��8O>�KgܐįCI\����������UmJ���޻�^�7�����8!�]i�1&��W�=����1,
�$�@zbmNߝ�L��˭&�Y�z��- �X�p���䟝��䜝���cߊ��Q�hk����X	n
����Ò�*��v����B�i���;Ģ&��E�֢Qp�D��D��-������j�F������a��/J������@�<V#��EIl��o��hޚ;N�h�"��៳B���ԟ~V*�#��"6h�g����I[�N����ԧ@N���ѿ���efG�I�dq���i�����WH���.*�S�BAҭq��/����/s��^�Ѝ�	�(��o(��/n���NƢ�I���?x�z�hV�/�y	���7��v��	W�% [�AQ�)!�ݨ`�1][+��@h:��M��=����X*��^m�
#����#�*/$�ގ�-O&��s�u=��Qݘ˺�W�x ���g-�#�^-̈́'CcW=�{3�%Ҁ��N�W�\���H�4�9�2���kgv��5�u�,�֡|Nc��mh��.0�M^B�D&GXG* ���>e�5+�q 41B�p��J�� �L/}�X�I����䥸'���2>΀Ka'���snG�����껠G̗tڊ'���L��}��/��L�2���7�I4�n���ڢn�h'�6[�J.٢��vƹˈꩾ���n�r1��(PE�����9��S$t��]�&\�˻��O2Xp��k�AWp:��DO���`�=e[�)��]��ar� Q(��.=��}]����&��{���c��9�F����hw��n��� �"Y�6��&J�7�"e�Gz�Ǩ�>���J{�p����fZOaYb+.+*��Cl�o\}Ŭ�B�R>�%J}C��|���]Z�[�m��K��ݚ�EKE��/׌"�,��^�H�qϬ ����b��K�,WGɩB�0'��]�멠ܗ�l?p�)��Dj�A]G��X��`d���[�����gr��M����ǵ3���ȁ6Y�]M9���	�YػU�6�xK�m:T��Q�=V#�-�#X\p+�YSVn�L}���E�Ht������=S�1��2�}��ˊ��%�B�b#pQ������:Z���C%(�>����q߯	����~t�E���
J�{
�3u�Eo���V�dK��e:�Q[�.OR�B�D���_#�j�T^�D�P, �n(��l��HI�$T)Y�itMy���я�x�7҇o��5�C{��Z���Q?j�)L���"�=�M ���lq�G��6�l8űH#�zx9�Av�%�r�Hdט4T�����_���}�!��+��A�z�Tn-�S�^r�z�����O�H����	�b��R����E�g��V0G����C|#����V���yip����)�9�kѽ�Ċ�Z{t�b��В6#w4�O��ݫ�^^e�K/b��V�SiO���L�j�R3 A��.���p�	���$���� ���$c�@��7���.b"oW���o���4�sͬ�/M��
2���>;N7��W@kO�uB�Cυ���y�b��\4�	�D��{y�����7��J�4w�X�M���J�t�$yO�%�
t:��tC�������X��N�~�<���p&�	��R��1S֬���(����He@�ӄ���ed8і���Ù��f�D[5��T�)�g���"��	��4��*��aqI ���&Ur�JO��Z����ƿ��B�X������z.Rx� c��c
�6i����O[<ȹ�����~I�b�
 q(�d�J��o|#��=Ӏ�)F��+\
�(Z	>����i���wn��=4���9B�(u����)��I�`=6��xq&W�Kg���5TR� -����i%/-�C���yR��98-����)F�Q���L|����^|8��2q�gB�kw�>J����jRCF��MA�x��D!Kn��Rݙ���llk����1==�5,�P2�;90�y����NO9�d"�����/kb/(����������[�fx'�%�ѯyf4��^�q/�s�\��o�=P�����TRϔ�Z�r伩xy�����NtS�@K�D���Zy;�s�����j�짦��wΎ�R�9<��U%�)�beJy����w$��К|�	2�<r#�M�C� KBh���l�PݷS�ma�穝�F��-���̪���Ⱦ/���q]*��#"���)2���W���5)�����]��p������IH��������76� F�=����#�7Ԛ*��˼�Q�5���_�>�;@SQr5��!n�*^י���1�ŇO\�~�$���oU�/N+~�
��`�ȡ���/N@�!��|eg��{�nl�7[��<��#q�������ѡ$��Kr�$�LaQ9�������^��[�������yf�՜ ��������-���DZע@�
I��h�4�zf��2�GР�C��h재A�vA]����V���Z�����,��$�X3����;PMiD����X��{Ddb�������j���7����q@���-�+1��<��#���"����V��"̄0�- ���F�#M-O�ʉv`���V������C�`��>t�;Y�O%��׬�[�Xϊ��W7�Y��NU0f��Gq���柿�|��N�	y��Z.���)�yA 
�A��4?��/ѽ=e�|��4fI��듉g�Ue'P����-��F.��K���*����k��r"�N���I*ި|2Z��(8��Q���H(H���{+��,s���U��Lz�i�ţ��5e��g��3�������)��Bi��;c���8(��b�ܚxy�do�W��5�X�&U���C%��ȼ���u%T*����C�{�:Z^������yG�jX�D��W؈Ĥy��F�C�������F�"��Z�M�,B�b��"H(��J|�F"HhO�QtY}�>��0;�ޛ Jw-�ۓF�%��>m�3��������;�I6�O՛5�_P��82��'�aNP��T�5���)t��?j�~��p:��:����#C>(�M!}[<�g����F��I����&ȗfUB���;G������j{!;,��v�ܸ��J� $6C�Z:����J�p�߫�����ȕ�]�s�>���u��BT-�Qz?����	�VNҠ��}����������%_9�t�RC�+O�v_P�1ϴv��vb���É-D9��d��e�iF�t���D	�4��R�_$��~����0�b��\f#��؎�t���3S���]n ���5���-gtm\>��.N
��1T��4�}��6R��m-��� �V �#=2�'�p�?"��jt���~��ƭ�#>+m�nS��#}x����Z,�1��v�}بJ�#h(�*���b��Li�Z��I��e�M�ni(-O"��( >��ݱZ��iX����С���i-��9R��.&����10��ǘ�2E�b�_���dDt8�N�-���u�r�J�i�5P{����'B���U~��
O����R���j��#|�-n�z3%�a��hp��g:`Ff��U��{if��P-�0���0�� O�Ƌ�f����S�ր Bه�,s�{	�����k�T�'Zx�.z�4x����u�r� ��Q;*���'��+9B��I'�8Ԝ����`Xܖ�?�p��ܿи�ԖB%7�ךA��C
zSښ�ł U�Pd6���S)K�f��ZA�_fp:\��~��6��M��矣�O|�t��ͥo~[)R�jG���B2�%:���m�shp���l���D�������l=\�wͩ7��,��5:�f9�Kj��.9�)�#����ʊ��TNLl
ۣ`4��nR���|����@�/J����3O� �or��kꈦ���OV��k�UO��/����ߕ_���___����j�Lh��=������"t:{��ba�{�j[
�6��r�H���ҵ>�Hp-{�����aJ���s�����ͻ��J�q�@ � *�'��L��,+h���~��H�R����6�]�����+������r�� ;�<��E.�$�Ϲ ����'־4��h<�<ï1� u�mN�SZk�k����t�6���e���S}���飊��$(�h���Y3��<U�A�5�cku0ė]�5�ccC���)�	S{��)�]M*_��SU��a�J/$4d�������]�a�k��e�����=-.�#�@@��0��AN�,R�ԋ��~�S)7j5σQ�5s�Gx0��(��q��p�����͘�@�ϫ���)�����7��{����@�Yȫ�PB+�1cM�\TH]>��ſ�F�A
�)ӭv$.��4$�Y���M��D�����ү}�̄)������T1H��f4������w�~�6No�x.o���~~p��l>����#V��&"�/�ܟ^:P��gu�i���o�w9꓄R�{.�"������6�"M��J ��oX������L�d5���8\c~Ú���w����6��|+^��,PP�4ډ�������b��*DK;�>|��a��ڿ�Q([���~��]�ͣ��Ei|���1O��H>�4) �TXD���^�Ÿk�R��e�	�{�bI/}l�a4��R�t�'��Aj�2��`^c��[���>���/$�u�}�?͕a�d�-
d�5�ԅ|�vէUv8�FO�=�e�ˤ6�a����2Pw��w*���.��4:�!*sAf��VY^U~����Al)Tf_�����IH�C��	�d}�{b5�d�|�B�u��ys��H;0�����$���VD\n9���5�ݠ�y�,���X�9|=���~&�KƏ���U��} ��ͭ�����r��$&�I��FT�?n8o�H��Zo�Gk��&\�g:�;:�v���a�Ic�e�g+{`����,�j#hE��I�a(t2 "�)�٬Y-��R ���p5��22���gJ]D�|i�
Z��)�Na��;��l��JN:��Ý�Ny��;�5:mXɇ����kҶ�u�ll���uFH�j0@B��;����=���U.d_>Q�>�,#�����u8��of��`nD#�J�UX^����\o�3�[�}�U���ņ7�6���mE���'��Y��@�Un3���Sع�,&&�C��p�5��P�(M!��KO��7��?k���~6{�+��|O���7�xڷ�ph�b�э0@� h�p}?��!�m:)�~�4��C�z���U��13 �f2e��8y�*\e?��@���*�3����Ԑj�J��$S����4ʨ�a{Ǯ�H �A`������(��q@Gz��zX ���O��-\���`I.�D���]�Z��r�yg�EWt�ݓ`��6��P�y���ϚeEb��ʑ�ο3*Yp{/`;������Q�[*9 ؟��0y��2����Z��s�cm ּ?����aG�dk�ɓ�����%�(��ɐ�Gz7CmFa�'k[`T^�͠��P6,z��,E�=�-���B���Bڇ�|*�(�f�ʿg�c���Cl���Ds�,JM7^�5�-Ηp�<���x�i���u{8T�8��{��b������F}��~�E�-Z���5]:Z�L��j3��aFk��G7I��ռ��>]�bS�#��z�!��ZO��L~JM�j�w��������ܻY��0��IpEw���FȊⱮU��̛�)��Ǔ��-���|��ӯ���;�;��	۶y�ĕss��zh��L�0!��=pW���W~f��P ���v6��	���Z���0�̗F0>�ƨ'ZpI�沕���d�:]�_.SI[��[=j�s ��@�9&��L`D�"q{=T���5�D�����P��M&}�c$g;�' s{Η�*��)}�x�q��]��^���y 
ɗD'}���q��G�\6ZhK��a6�'��v��~�$A��b{ �`��؏�&����u�嵌�K}щ���7��ۣV� �<�o�c��쬾��0��Z��Y�����f&?{uD����1�1�}yM��{%z2�:ǳC�9TJ�	���[�&�
C>�2u�~��k$�:j:�k���E��]����Υ��_!��}�V�v!�Zr	0�d��M�X�Ơ\C����[�S�FB�'ctd���_�E$���8I�n�tMI�@8���H~��<ޟ�:�<1�?�tR���^�ͻ�;����ά��N��3��G�UO��sd15uנ�q���;���|>�k��Z_`����q������?��ǖ�_n�s s���3���K;��:��mG�&\��0�aSZ�{���J��+���X0bEb?޹���G�4~`^�&�g�(���q�=�_%BO.�ה�x�����&�#�'��o�Ӕ��d���&�?
Q�q�+�ʭýc������,c{�nK��g ���k���t�LŹ\V��Y�)���<��{}�h�yi�絵�� �9aMD�����k�4��}�k���y��F��`Đ�K�ͫG �����q��+�z.Da���Û�Q�:>=Ŏ�K�Y���s}��7�&G��'��/�^����(�etsaq���ﲄ!d�+l&K����ϐa��;�$ ��d����ۑ��֑L�(���c�ר��l�c"6P�����2�5��e��@v�w�(}��7�Z�5X��ܶ���gL_����N���K�+�Ɨ��#M��_>�xs.�7�O	��6���[�ߑ�p�<����2��И��q����%e��Xɸ���w{n7����ժ��&�����3����J�������_��:ME�⊚�g�����D{��R��DT��:��o)�7�X�a�;v��k7Z��r�>�J�hDH[������!��$?ݮ�Wn�r���z�6�I87mWρޣ� 4�\F;L�V�����N��Y�dezMK2G�����5w���׽�,�.*C>\� d�w��0�Yi׽1F���r��;�����!���,Bq���O�
)J4Y��j��]V�:Ivd���AZ7sȀ���^E_�@o�6h �W�1O�/��iGN�e�>)�=��%?���<��E6���J�I�G�N������Wv�;f�SCョ�&3���\5�o���[�G��G�g��L̫�mAFT}��Q��_�!����g�1���m��۠F$�(N��?�;��8;��b@SG��?Qr�A�ҔU+�&�6��͜����%�/ʞ�Z�����	�i��	2(z\R�a]o$�!�!tC|.*~�`�䟯���.��1
�A8�٦ȠD1T�Oh�7���>��彏���C��\��2r�����@Q�,�������G,�1č)F���5�d����5��:xKeQh����ZZ�6ś�Y�5��@l�{$U��0�]u��1J� �DP�X7T�_��yT��z�81fGď�NE� O�\菲X!��.~�l��H��Yb��L�gN��|���T�J [��; �b��Fm���\���?M�B�-��\_W����b���%r�v����.�n^b��e�_��{ȹ
��
Gx�J��i��0-2� �۽��U11���(�)�(K��n�S�C�s{��9ZḴ1�㹖��JV?ㆲL�2@�<sOS���l���y�:���y�}Fc7��Odtwc����$
51��s?�=�k^�k�S�|�@D��'z�݇�Y(i�������>M��&�=���,�}-��ϖ#ʌ�iʃF�0=~\�ӛgo}��gv��GV�o/�(W��__��ĺ6d%��"�,�-�mx^&*Q�0��ѲpZs�[1�Y&��}/?TL"��M*�j>��� ��H[�o���]�6�5��̜�F᥃��R9���Bd⟏�[��ƚ6�y�ԫ�GGsy_s$���:���� ��N�y�"u�UԶ���G�v�T_~�|-�����1\��c�r/;}��m�)�b�$τd�^9L��1��h�[�Hl�5��Hy�jZ��~��8��f\2n�_�.`F���/V�Fg͙} h�h��O�t�*�V[yv��\�-�s�`/�Ƥ�9oI��4FL2H�qf��R#>�>&ftM��Xi���D��˖���Ax"�Dߠ:'t}^hMiqP���Y߯�����o���L'��?�09l�zvD�F���{n�?R��u�Ȳ]��дlmD�o�܊y��g:�;u�slDЯ��@R�XG���.�!�~R[��W�n�=��	#Ed?��O����o���h����Vz�\�b������)N��}��a�_Mz��^�U�2ѽ�Z5E[B�AKwhݽ�ԯ�?�5Y��AȄB��2ϯLkHu ��>��d�9S��v$s�?�GL������Am�еJwt�3��]k��A�ԋo�P�ji�of���Gk6F^�f?���$ɏ��P܍�P��i�^=E����m#1�ҧ�N���z7���&�����f��o}���������L�>◱1�w�j���7����^H���O܌��~]g���T��")ce�K��x��2,���,��elZ�ޗ�����S/됹f�c�,>(Go�`�Ax)�:���G{����̪�$��mO���9�1��Є�7I��@�vR"��Ƈ�C˨��Z ©,�o���Rm��_���1�V�����8�;������� ��~9x���&��f��f$�A�WG��jm�:�����..	�1�-���"<����'i9�%>��	�5`� ���+����Γ������O&�Ř��# ��C3�M��uC!�Cc*e�q�jⶴ���{=�w��)#$$}�c+^ ��S��?j�;m�XF�2|���6I�^�13g��.D,d;��+"�/��T�;��܍�4�[����^;�mE�9m��~K��܆ѿv�؈���'�Q��E�bf�n+e���̾`�¥�s������x��7z��@A���r��2�N)q!��
��[�� �{k�t �}c>�5>nBȋ_6��{��.mc�X�<��R��b&o�����q3��!G������_��L����g��A`��e#�@�Zz����T,��Ix*I��,NR�5.��� Q�,�$���g�Yeh�۲�/%���7
B�p�0�?z�& ������V�G���n�}��F���O�wڼ�p���V���ؙsBR�=��kI�=��k�e_}
ؙ`��g@��FބŚ�l�ܳ[W�q-�E���w���LP}��Eq���x��r\q�E��$�#�6�� �y7�ӿl��~v���R��`v��U4`��[T�޽̼���Wt�mp����1�ɫ���G*�ֱ/�I.���Ժ�U�RO�m�c�]!gRm�6��LK�����l�߀;�0 6�>r:����8�N��<�W�U��7��m��n��ѓv� ����Bi,(:cʹ7A�~l}l)�&1e�{�G�
o	��������z���˲�,� r�N&�h�����dZ�43�Vh気-��|�0_h\,cp�ab�E��-Ԋo�[C���KP���������4�׿R��D�47��Z�D�������c%�ˌP5����4dY�13Nd���mV����c���n\�����}7����*�|;��Z��خٳhL�Ng��|�uk�Gj`jj�o��
G�A_t�$w:_��$��%���i�=���U�rS���5ȉ���N�;fPX��@��W>������
�Z��0�6�G��RUp��1Ml	�R��(��d]����~l v�M���e�é�.ېp��[�r�{���V�^bC'����s�)��N�b�dԣ��ΗԎ�D��
��M��T<.|6Y��!&�?��(F+f�u����������0�~}���Yܘq]Z���s2�D�5� �I�XHT�Ԍ��
C��k5���@� o��QЯ�l���%���&�eJ$"H��Ѕ(P��J^�n�;#*xGE�+���طHߐw�|����ǏN�14,x�n�@�o.|��wpt��,L}h�-3�N�0����M�{�VW�.����f��l��K�#J[ă㷂�+�m�h��7;	�v]�C�no��n;�mdMY���J?��p=�S�"��t�Rs�
�|0K�d��=A�,���"�=/��%n;YGn�y�FL��J��6Wn�o��
��l�/M�쩑���:�=����J��j�F�9�4H( �]��PJ�C��n��C@@��A����Cw~��{���}���+f�5�k���7�cG%�,ލ������=mة�B�d�\淘�;J��`<`�H�qEP�>���� 8D>,�}��]��3�@pB����*�������w�T5����W<�Wn%<܊[��S��T�+q�B�	YKM�X��v��j����qO���iu��܏Ƕ�����âً���e6�����ߌ�h	(3�5�� :��b��nf������ ������Ñ_i�������I`��'���L��"�n	�t.�K�X`��ۖ�q��_y%�9L<�7��ӑ���?(����з���>�6����n��俎R��s�w���&�M�~P�L��&�#�+Ȣ�aJ:^ݏ�ٜ��b1�I2������W�����R��V-�V�s�5�hyq\3��?f=ZG/~�ۺ�ȀО���<?G���6й��b@D��8�F�65�y�C�jcߚ̓"���E�*�qy��!������1����~�'b������0���Y"��w�u��`Ƶ@(��J;�_�m�d�{ך��h��PU�{�q��5�?��~��+��M 
��e�~`�·f8���0X,����8�lo�w̟�PG0�]�H�����w¬P��Χq|�{uS��"6ETxP�1?�^,�(�w<<�[��}�
ͥ�XOXLu�]Cc6����8K+ٱy�!s����
����C��կ �||��ڼls$I��+��%�C���I�is��{=�4[�m�O` �)~AL
�xnִ���L���o�K*�!�l���{���3�/����V�<�_G�����/N�*e�b�a/�*�F���%Ӻ}C��Ȍ�ݬ�u�(c:> (�H'�o�~�s)�(J��c�^�/?v�h8�E�����aNW�_�n]a��%�T��-�����H[�s�қ'�,��l|�a"��à��\\�Tg/M����'�P��ص�]�n�y�lG딑K�1Z]I.Ѹp.�M���v��[���W��9�~��8-^1��0�M��F�z��7Wi�W?����m��8�!�\h�/ ��Qm�KRh8[)z��nixק� h��<�{��e���7\��H�ΎDf����I�v~#��n��4�ϱ5�����P~ebk9$�3����%L��BX��LZF�16 	A��+O0z�~���FǴ:t|�}�����ԑ+'	y�}B^L�� bNK��v��7��d�8��Y�z�@1y>	颉�����|Z_�hK�g�!�<��}Q����3�5�$�"݀���`�Sb؝GW�m��˽4Ƹ-�~G/��ϵ;u'����};P�e�� �o#�6ͩ,�%����ܬ�a���u¢#�^C�׈�#ךVeM��,���$X9�q�mf��%?SO�}Ej*:G�[>�y�	��Z���b�Љ��ػ�E6E�b�� �ה��������@��@y�l��C�hw72�x��9K����`�`��8�m����l24Z B|V-<��7	���/r)��0�{��x���5M ��F�:���jV�F����I���H�P��{�����x~��غ��2��vfH�tOe��f���yfHD��9C��)5� ��c�9Ŷ�� �1sB[���$��1��JA��ۏ�:��):�*�O�O[b3���i_jZ�&�Ǧ_�t:� �E��~l�ا��`�G�5�c<�k����$��n�bԋ����B����NFغnm�^I��M�z�_(��� ug������I��Pr�x�&�S�u@ �N�Z���ޙ���7��l�xJ�P�,��y��4�8w�o�P4#����k��!�5ٽv4��6��������.�c
��h5$�����(�hh'�_�4�����S����؏WW�\f	�
UP['T�-��f�bI{�~}X!H�<D�w__�ؐ${	Hil(0���
��0�g���a�4"h�����r�3��t'VM��"s�5���y�Gx��5��p9�qYy���
�=���)�� _�&�w\V�m���wO��U�O¯I#�F5�����-8�KE�.�z��M��Ri>�ҷ�����:_L��(K�Y뙽�M���0���ȧ&2�	�X-:��S���Z�P���f7n)JK��������[�z|�-Q3���&����È�A�*�_�*nM$��F�)��H��O�bk�9?���$Rg�^�Ժ��}�_�:�9���΁���.�Z��y���,�窩*ʺ��YKLa��b!����$���C^w竽�eu�i�����o9t�W_vu�^T���\H"�  �,w��֓�Ј8�r�%��.e]�,��J�2���Y�%g�8v�Zn�;Ȍz75k�xI6����91e�ܟ[-SH�D����p�Bb�I�ǼF��a,��9�E\�:��&:]�A�#���;U�D��-K�il����vET�r�5��us\��;Qͧ7��f9;uv�^Xs����6�::PPj_u��M��'UͲ,V��~F3��V������S'��}�v��{�4���i�5����X*1ɚ�B�G����#�������qi;u�HUM��N�ܘl�`E�/�QX����.�d�<}�	�%\g)�?�f�C@�wD�n���b��"���F�����EíYa~�6A�c�Qj�S��#8��1��[�0���Y�Ay{E�cn��+�*�mL��L�@����C4�ԉ��o�3	
1��R�,�M����&��:��H}�ܿ�o�'i�?�Z�r�����i�j�
`j5���C�S�n���~x�}�/�G6f�3#(��~993 cqr^CNl��x}�$�m(�3�O��x6�jzY�H_'~�W�R�W�y�C8��F���8і�R+%�;+R_�W4�h���r�S�|��HIߥs�}�س���Su�	��[�x�������a1�s�\�\n����֭����>cG�_�>��ld�
ƜVҨP������B=vp'e|�l�����@և5_�&I�7�L�LuNo��褼;�R��*D�Y���c��b�!'�,�£0qV|;�U)�W��5��ٷ@�}���n����Xr(z�׶�F�ʣ��l�a���ŷW�Ҋ��w���W���U��J�K��M�."%}�*�:��Vĵ�E]����6s<�v�.?�\��L���W<�Wg!�����R���2�6��6��ɗ����L�V۶R�����*�r�j�Ӆ�њ��,��&t7]{-���;�o��j�����9��0nu�4f�o'��{7��<P8��H?U�I�I�ٿ.(h��L]1�$�sH��v��U���߷_��X8VS��7=�.:��+��j�IJ�Q��X�����5v)#�u+W�i1�q})�['�/�s�t#�/x����� u���tWT:��VE����W�*{��p�I�O^x>�|��v�ӫ���ŒkԊ�鉌�mUj�����Ar�m���9�+��`"���rxѾvЩ�3U��y��&$}/�Ӯ�c\����*o/|M�D�D�[��H�!7N�Y��$~�s([K���òu�کB<�}Y�d���gjN�uό�v���U`�D�ȏ�Ϭ��6�WR�s�^����O_(e*���X�����u�B�5^Km���C�$<'�S�u�S�h_t���.pmo�j���_��(J�LPI�[��,W�jq�k��Y�!]?;rd!LY��r6ay�ة���~/������q��p�Ke��j���n�I�ݜ�Zǋ�h���]ƾ�ǧ�KZ<5mfx3f�Tn����w)y�v��h��v3ł_Ҩ/���{J���7?eg�}G�C5f���TF���4�0�4I��_��Z]� $Mi�b���-7:D�ִVejk��Eu\_术�,y�itwJ�+�u��Q�݆|)����F/�5?4ke��v�3�Ū�"����՟���^�K�I����m� �eY~�Y�g?��i���ӝďP�U�c�57�}�� N��7V�VeNL-SpÁJs|�[>�@^I��M��4�2Hy`ro@�s&�X "W0.đ#�s��I&�B�!�E�g�%��$�{m(�/����� ��<�A��4?8��v��ЭI��28Az*S�=Er6�1�_�7^�K�U���~��ÄK��v�S.��6�����u��oHQ@�v���@>�:�r皴Pm%� 84)��8$0ѿ���-ͱ+#fY�p�{����Ԡ_U����*��T����XV���zTt�z�C�^L�.�On΂�?�s�S��.!UO�49���9�&����Q�7���Ӈ��B�yi�.�Hi1Jn�f��g_����1���!��`J>f^�]��~@�Rn55%	�L��7i�1�kqy�Yȅ]��	[g�/�a�$j���*s+�4�_�n�w��Yj 㬇�y[*��V�1�����$˥�5zg�Ani���\��B3\y�P��k '��u7<�ϭt����f�ر��6�!���&D8~uzU�\����1b�w{���2��v�¸�xi'�1<��J�&��C��׷.Yt�epꙟT��k��Z�"m@tB���^p���$����*;bNP�=���l\����g|��������G����'M=����R�Z��'�\�������D�cL��3��i��c�ҍ�	uٙ��䫵����Ra`�E�T-b�������#��T��ӽ�"8��S7�R>�ju�-�f�҄ɀ��y�"�
���K����6?N>D���B��W���L�t�����<^t.���0�%pW>Ƨj|���M�+?�.�H��<y�Q��2�����>0]nb� Y�T�`j�N����}*�%vi�� 4����a㺐��G@N�46�;F��wM<�+���a*
E����ґ#{W*�$�+����u@1���,^É~���x�1�1�f����%纰q[y��<�=J<�S��]>���a�?���CY��ʌ�f7���FZ���P;tv{ts�1`��Ҹ��k�����u-g��yr0���>�w�k,B�*�p$ܣ�������kv���u��eb�}7�?�����c\dq��R����w�%O��P�
�ȝrީjJZ�
讀����3���Z����u}Ђ���b��N�i(�nM��qg�k�Žʎ�~pʱ]p��z�?��ߚ*ȶ�K�"�k>��f��V����ú�$�Q1��	��l+�%p�r��94��Y�4b)'b�8�BjL���#�.,Y��ڗ��f�}��\C��M��t֗��[Ҫ�X��Fe2��!��i��T�Z(y���;�����L�O�曋*�:x���L�_�Z8Zپ������y$���������{�_�nX�1����H�ԉc�
;��[7ő��M$����bz���>(����S��^r�>� �j-z׬Ȇ�s�n�
)�G"Q�.�=!�I�/�왊$��ᑙ�J�6_~��;�gV��oP-�U~}ʂ�+u�f���~L���c 3%5��4$��%��ݼSl;�I!F��b��Z>��zU~!	(�|�jI�j(�j���P�1���!h��j=�������Z�ʘ�g��R�F�'G�u��F0�;I�L��@չ'U��CC��e�!�_���P��#����U,Ƴ1�� X���TQ1�X����t������E}D9O� ���R�}R.EV���TSmս1��xP��j';w;�lwb�N�}��灢��?v�2��Ұy�Y��9��XI@<D0�2�2���Y.(��h�#X�X�J����ː���ۑi�g�)��J�6�Ixj��X��\��u� l��;���Je�n��+"���^B���n��<ܐl:Z9yB�p�a�EE�4��L�Ǳ�/>����gSQ.z`���{���f²n��K�i�Zr�0"�L�j���`�ئy��oA�(��v)�8�(�`���~�]�:x\ )� �D��>޲PY��驖b�����8���vl~�� �B���ۡA��5�|h��ZA&�tGV�O�G���yv��}���D��x�.�$��{��v/�ͫ~��T�3�ux�X�n:�{Fn�%zAO���4�>9ţ+Q�bq#�`xJ4O�2;�h��G�OF��,�ꖑ���8�,,9�E���Q�f�Nz����G��V�^.�R�	lBݖV���:vAn���&�Y�*�=��醃������ώ��oS)`��M��ڳ!��Z�e� %�?c$�S�7z�ׄ�����B��߾��B�
(�F����L�obt"0�2��q�`]	yP�$е����Jܨ�(���]�q��{J�� �"Sǁ� ��&А���ЈF%��F�w6='^n>ԎI�%�x�K��^~�|�[1<T�LOu˿	�ʁ�;`��[�ތ?��
,s�]�	�{t�ʿ#F��O�FH`��� �@��W�S����pL0�<H0�EX5���V�?�Y�B�/�� 뀉2Ҁ��x�	��FӉn�.p&�U@�L�7�-�������(��1���9��`1���7�K� {=�V��VlA���V�VPaA핃X����|� ��	
�l\hh� ���}	J ���Ue��J��Sy��|����oĹ�C"��w=�D�ƍbq*�[	�-��]>/>�Jŷ�ߵ��	BU������z�m\�c$��5�"VrLM��U?� z��q��e�J���nٰ��7R�.�/�=<9\�A��8F�z�������Kf�	� ,��L�S�٠���vtJ���"N��ޮ`[�P��@�Ϩ:���[���ި�u��t?�P)�bTt�Nަ���w��=^wȮS���6\x�9�t�����D��"����ay�;���@�qH�����J��C�C�?)��,����8U�ğA���csb�);�X�zMΏ�`ĕzpkР�c��	<I����M^��!���@��|:ՌY?L-��C�8>�U�����?�5E3{���ly|OI,	��� �/�=(f����Cw4��Oy������Q�0N���m�˅�Z}#e[��-�GD$����PG7�� O��S��D��0J���b1CD������aVbf�>"A����cT!!˄H���E�S��n�Yp�l*�W�NIcX�f�k�Bme^�N�A����q�s��R6V��x�:��q6��#@L�`6R��]�`�z#��]y�z��!���u��%���,p���
q�EOCZ��^" �4����S�"o~�D�2��m�%�3忔C�|�X��� �Q���Ċ�2��!���6V$`<��:U,����B�n�Vшu*�j�k	w>��:��.xL$v-Q��w�5%� �ᴀ��7�T��p�����8�Z)��?�EU2�:�j�*R�g�wx2��j,ԣ�]�EhAO����!k8(�f�����)EH�k=3�i*��[�/�L3����𫭭��N9-���፤�u�D�9�+��P��'�"R4�e����*�����ƿT�"DE�N�����$Kk�	��UoE�'?�,��6�)�ȚG�>,|BCޗ�U:�pvX���V��
'�"31Yk���2�!�D���o�>pN�?��n|���}��K���O�_������]$,pIP��Tp ��O�T֔���߆�k��)b��S<���o�wCY6%�̢�if�ƹ�`��|�����J�5�>j
/�m̊LO0��z��\�U�o�#�G��p�b�"�&��!�1+Lu	�c�[�ύl%7�L��e�4:1TDʐ^PF�?���q@�}i�uok�veD�'��A�+� ��˿E]"?e&�-�Ϛ�ݻ|EO@]=�MC�=�Ԕ/�j/�����Ν�J�u��A{%z�)��,j&��B�"���2�+�	�"&�m�������Q"�$�d�(�p���"��'*ھyk��9/��&�IO�ޔ�hv��OV�kQ��Ax-(Ti+��M��FK����&��c���hL��N0���[;�=̨�#�����f��M��0n��kr)Ƞ������ ��{����!o"J�`�[֧�Q� �9BDt�??�����܏�ɡs[��2vs�}���O�p})3����{�)�o(`�_|Ǳ�����8�'�5����,��_ɔi�b��ZZ�O�V�����QTm>	~qINާ�� ���v��:������4:O)�f���޹��;��r���};Y!�ZN���B�2/|��)���W�IyA�'�h�au煎mGqxs)�3��Ѣ�UH�jjZl���+>��6��KQ� j�,i�(j蹊J(�X�/Q����������cv1�0�?���x����t�ȳNMmmk	��Z�|  �&��@�V`�T�j�������l�������H�5
.��uk�f������n^��wKNWc\t��U����*��V �p��ٍ��ڭ~��#g�cr=�T�_�c�D�ظ� �,���D3[67S�A6�6�|>�`�kF�.ǳ��jd�ae���y�分f<cG�egF�ܶ65ި"8,s_���m��5�*��\�\8��D�;0D*��`�U`�[�F��O	�m�t>!�Hn������o�]k�!]�^5��W�w���H0\�:#��eu]p�k� y�J��OМp�5Z�_���W�#�tY��:W�U���MmD��:��J� H�	4+���f�b�Ģ���7]Z,?j��T@m!֡�[{)�u�p�K���?�mz��i1��;1�F�����<�񢏭'�z�jos�[���J2���n�g�;o��r�*ì���H�+R�.P�Dg�Kn��(�\~�,�w�����"�Vݬ������2y�ȧ`����(���.��R�>`�f��	���s�{�{�v���V�.���Ϙ��6$��ma\5�����^�_ 7�$+F+
��U(o�(*z�X�^���O�d��K���x&%�S�<�l�z���DcO��A���Sڵ�pCvu�9C����z;&�����k��c���6a^v5K�������n��Y-j�=�B�T������۷ˎ$�����NF�>t6��YnYx��<�EQ��9��]�`��'�Ǧ�3����g��ݨ0$nv�H�Ӆ� �����Y�����O+��c����F��C���z-�k�_�6������GXҁ��n7A���9��?W�$	�������7ȳ�UM(p���Q�SļzZ��
��&;�P51�T���ɨ�� x�ۏ_�d�J9�!��a�$xgX�q��O��h���ѱJ�{R���N� +��2���)���ҹD��G���:�P����Ѩ����z�A���˷/����8&d����z�3M�a�vԿ��@2�W�B��1Ղ�(E�# �X_�K��f.�4w��������
	� �[�~U�G��Q�=�ឤ��E?[0y�k�W�U'*5���^���*���ҋ/�Y.K���~���`t�O�6��$��We&�tnbub��3����*��1�K6)7o��ҙg�Q��+ڎ����c�1X,����z�q�_��?�a^<�8�^O�'w�Aɢ��Z��h[���I�ؠ�}�E�&ki��ܳf�2�a��˧�5�S߽��N��"����R�����yTwZJ�_�}�=�$YɼA Fn���C[|	�5>�����:���-; h��%����47��(&h?N�1�����yE�~o-��Ř�>�Zˮݯ��N@�1��R0��l��\H��
�4���X�\�B'���+֧�^�ǿ��B�q�w|v��rkMg�I���#�xX�/��Ǽx����ɥ��p~�'�� -�����f�����L�:������[�{�湰CC�m��i\k�t;-|HCN%Mm`q�&��=*���j�w^'E��D_!��e_$g?���$y'��3�5�D�"��A��II��3s�T4<`�G��!�>�������1,���~����ԙ��w���;M�}͟�z�9,�=s��|̛�&@CboxOb�wC}=o�`�D��́�}���Z�����T���{W�
<Vt=�G����4�ba�^�B6k�'w(�CS!�l� �V�k�� L���ʞ���i�|�HCV���XkY잍|�,��@^��.�'Q_S��+bD�z`\��-�/
:�t^����Y���:���RUt��3��6�q��A���+=l��/T,h�9��ĭخƷ	fԪ���c����ε�H]kh�8ϥ�:�WV��ez�.�'�$q����R-@o�%�J+�}!�E�Y�`g}nv,v��y�]�&1h���0������ڧ�&�V��sZձ�&��G��*tº���u�����|GR6�������=��S�O/������Tpmð,>���_��Hb!��ݞ�%BšX�W͵���s�2�o��^]~��l&~k�^�=���p;�z�Wp�Ǵ�����%>�eO�[�`�?rx#�����v4�PF ��w��QS� o�Ȼ���d��Q�:�^�S����A�q�<<@^�F��PP��l9͚v�U�z��5�'�>��g��.wX��A\�����򓑾����Y�Vr���z�aI풮��8�%�����C��z��csQ m���a�]�^��wC��|����/�:�s�4�vTE��:H�Z]DՑ���`H
صhOGf-#�DI�5];H�T��H֚� ����4��8P{�d�d�Z���doO]���$��u��l<\��}���߁U����ο��4]��ŅFn,���N��8xCS?�1w�:5%%QYj������D���&K�n�4�[�j^��h��l%�ڳ�j#KĎ`n�ԧ��.q��+��*>%�{��CDnaHg�ߥ�b�n�ƨ]����&
O��
7>ϼle�Wld�Ŀ*�?�
����17�P�=A�m��wd�F(/2��sG�6U������i�U/�It�j�Z����d�Ep�]�+�����ӀZ��L�?�@T�L.-�� xV��M}��篲��O�"���\��v�O�X粩Jl�5h��k�BY�ݓ0�K����7�I��ǍȚ�UI�;��O�<$���9�Ɏ[2 ��s���C����>��KFB,Aц]F^A��h�.�1���y`�C�O�Fa�%=�+Lo �~�͇�����k���a_/?H�	��Q�c&��#@P޻z�^n�4�s"���IՇ�]��m��{X�"Hb`E�n�njS�9���JR0l^i���X��c����1U�Q(���9�@�;����@����<K�!'�{$���-p��Z� ���}� ��۹M��]O�
�c)��wm��S�ĺ�|��0�ݞ�(Ύ��(}�N����:b�q+��n6=�k��p�4��5���7�<+:)��$���b�R�Y�|�V���Λ��g&�m�קJ�.��F?J �K(��e���78UAw�6�w`�ŶO��7+aO?�Z��GH���q�=���� Mލ�6ج�s;)q��"����k2C�V=* S�0���-�x�b�� ������T���!!?'~�a`@D�'�<��b�fQ/V��:R�~!UC#u�����5�} �(���)�ZY�99]��@�g���^_[�v�ВK?��B{?�i�*@!���<\c%o)ʔ}j��i'6�a�.z�L�������|��$��u��p�*���XM�_�&K�4��z��&��@[�Ԅ=�z�����ߵ��@�.���]�6�7�pO]���i�'�']O{�u�^�}��e��x-5��"�:db��\�/�h	�gD��h"�"�~��n����;T��\a=��uHEc�x�2/�R'ų��P�/߾�ò��h��g�jl�&ވ'��P��<�@�I�n���!u��R��L���V!i���tMA��C�ŬpM^��׺�c�L���H|f��u�D1P������=m
�$�w'�B~G���V�f>(����mq�j����A�2!'�S'ǭ��+OQ���g~�.��^�Ԝ\y�{���N��6ke�J�T��\<Q���� h�-r�ċ`�<̅&���0b�v���r���}6T���N�@�.�j՜�Zv+� � )"�g]T������k��r(Q����T4�e1s�U���*�=���m�E��"����l7]�M��l�j�W���k�w�ev����m�о�i(�u͓�f+�R�]8u�)s�G[�fu9S+����T"+��̂�s���e�t�6���
F�%�spg�vU�/�n�r��7I�p�OQ��N
a���	=qj)	qmfJ��9�L�ǧ�����co� 3U��L�k�W�u�n=!��<��T�V���L*m�M��1�{�ƴ7*$��W��.{�s@�|�x�荣�1G��F�2��W�����A�Z<P��μ~q_SI�� �1󚘵َh���7�R����7=�qߞ�����+Υ�?�-4��5�z��vZ(��� �W�?>P�e�����3�MN-�k����oHGu�t�{˖��rq@/>b��ď���t�f�x�E��`)&~�HWy���ZN/n�Xz���7!	7���6/]Y����6� �lcN�)��DX�i^��ay�"���k�̫�^�K�>aO/�ޖ��aE��\�-�(�xo3��2����`(���ͅY}|��fX����% �^�Ò�ͅ�V�
�B˷�d���^�q�� �fG��<�X&k��,���	JJ��C��z�A�˫;n�-yy����Z) �b��f�ZJ���ڟ��F�_/�/��4�f�W�CPc�Fy�4$V�D��'���Fx�R��q��h��������ӽS�*�_��h���Z���������L�/;��wg4�چ�R{�<{���-_l�7�E�ǻP���\����p_��� 	AO�HND/����;�Q����>zII%�`��5�<�Yw�:�KW�2�#�q�do���jƱ5aIil�KЪ��~z��[�l��/B��ŐS����B���Z�͞��;&4TL��-OZ���Ȯ�Ȃ�pc©\[Sꚽ|��
Rf�Mk�/b��f���"Oq� ���ڵ
� �9(�`7D2�G0���r��G�2���� �ȗ�UO��v&2��y[��{�'�/Yx����^�#�Hy�-eZc�h�&-bԿ6�_>�_���H��C�]Ho��>LJ������
qbc��[�1��o�W[y��ú\��X��K��3���%k�->�;�*M�ŗ��0hR=|��< �#�A����ik�#�>�|���3�1~���jj�q�Qv�B�a�|��v�<O���K�3K)������
p�C_�� ϶���1��`���-V6!&�8r��~��Q�"�_XG�4K��¬QF�M^�[�I�����v�/�TUz�! S�Oc�$�X"	B�x>���3�$�f�HHc�Sd	��S�h�%�KI���mq�4e~���Ox؞��O9{WAyH쨋���G_Y�&p� �ȭ��N��6� J��`���,��Z�uqs�'v�cLj-��<"��w��'e�3�NV �YQ������B j�k~9�C+�7-_�8"B ��g�.K�|c�@�hkw�I�E�k99�Z�E�]JN��G�7���/$@%���a��R�.W���	,��\,����IT
 �
|�ŀ)���%OK��)T���Q�����O�٘���-WDF�AЋ�ӡ�o>=u�^����[��{����t��Y,w��V�ܺ8�q�%�p�s+�X.2oБ�A���D�w	���\����ΎD+��|[��������D�Q�@�%ɚ�����W�B�8x��іb��5��*A7�G\���߁X��4[|���@��:�^��/c���@�R��Z/��G�Ű�4�N�F��!�na
��;m^6�R�ɵ {��ha�k�J�*vO���:ʾ1A����,th ]�
��^v;�cZ�v?�?����
(���v�*��Փ�vK�'���.�&6��>������as�9�8�ʂ('�_#��}%�� 55
�쇡��1�`��2��&���7
�̺�'ۚU��S��[H��o�آN�I�:=o�����b��u�U��%R�c�����Y�7e�y�7J�+�L�ٳ#��7��Aׇ9�e'�X ӫ5���w��_kS��,.�<n������H�%[/N��u�K#�[��vgC*��0}�FՐ�����[�t�|�O������#�������h���ƭ9x�#7_��u��I�e<<�:��Y�@QT<U��:\i��~9����a���1�<��tx, �'
��fh�7t��+n�� BJ�������>N8�B��g!������h���F�x�5�������)a�����ɤ ���[�u�eg�@��b��c?	Ej2!�?_�2+/��[}6�Y���6.�k2�	]<i�̧{?��Sܝ�b��$
�R�
����\�jX[ݴF�����'�RY�{^���e3:�  O_/����������n+�產�j��Z�:�����g�z�PLE[�Q�j���|X�/Ϛ�?�X��5-I�Q$(tM��+���v$d��JG�,��ܲ���+��N���˴���oFxM'b��g��s������{��i��w��Q'��Q	ð4����n�W�/�L<c���0�n�W���W�c>W�\}�u�'�ʪ�}އ��?)<�%�G� �(��=lZ7Pȣb h��Fm���g�Ƌ$*���K�@&�vF�x�R|[v�<������t�&T��{N�숋3�(��Z̃���G��ar̎�]��㑽x��f�c~�Nf�u�����y�>�-�렓��t�)�P􀻽S��5�9��`��$�oO�AzmZ)&���+n��J⊓y���y$9٘�
3;�d m+C��6��M?;���b�?���@R�R�������G쟼N;�����,1��)����td�Q_4���>d��a�?�nG�{�ݣ��ݾv�����1V���<D �4�Y[�?6��$�kޝ`�w}-�7�GQ���q�����h�G,�k�d�bE����F���q۰�}RJy�r칓�q���X�L���R	���f���Yf%��rCvG�1���o!�o��w��Oc���ѵ�8]ڱ"�����K�[V������;;Q`w�X�*=���m�G�C�\��`2�.�#6����	ԩ���){�!x"U����2�ħ3'����&G��Z�xm�f����ט�8���_o�Ev��md'�^<�>�#�\�m
�# \4�<fD� �HO��e,�g'+���E����G�nQs#N�4���--%�m��Sp�.���о��͠@?.��<�����������g�|y �c��.�E��FSϹ��gҨ����Ei �W�c���j�j�"��e�wx�(]%,�	jt��RW0�چT�NQ�2F�mh�-��<���3�t->Ti��8vp#����@�BL��0		"f�Ѐ"&p�*�湽��u�O3�]ڄ�(��/nt-���;k��M�,��g�i����Hz��,�kq���C:���5�ٵ�c!�	'�p�/��Ā��=�`q��!de����j#�B�7���T<+;������iw`V-��"7|�G�����%�d��ni'w�"$�}��@��*�9B#��C_V��_�0�F����%�;�Z����p����?~�~�����ۻ@��ˇ]j�r�a��d��[3�ǖ��,??����h��8JTM�k��d�;������yx}��^f�uM����-Y'�z�tΉ&y˙���G�t��!�ǵ��nT���7z`,��m�lyr+�Jy}[�d���)~���ƞ�H����m`�z��rif�����n�N����t�ʖ� / ]���-�?j�3�#�0ӡ�[
5�ik�n��/!����Uz���S?P;y��q�VsB���p�Ψ	�\y�����pyP��x��b���f�Ԉ�a�H&�j߰A=�;�6n�Iv=��+U��y&א )+�{Y�+sK���4.��N^�rb��D*��@}@����kC���kل�L�ϣ$�`��\� �@c������C�yEkI}�B���Xv�њ�Qe,g(��F�*��#�SC�徎f�V-��87R���	n E�_��QW�4�Bw�o9�'uݗ;��lnj��`��(���M8^�
��"(Lk�8J�T�{{�b�M
)#cK�w�6��\����sz\��"$ �3���$W<S�#�=�|�N�%kH_{�a�� ��o�{n���1�m���GB��v_*)����Y�Mcf�o�79Ҥ'�vi	�r:�����4���Hӄ�М�"��W6L�uþ�<�1H@_d"�?�@�q�ٲs ̚g�j�C��i7��&�W��JW�`��1���J���ciue����ǩ����CيU�&����J��7[0�� �؎�,A�jӷ�o]Bp���XB=�3M'��q��i�k!�9�]�:Y#�>�������B��"X������8o1
~�}a��V�j��~r�*�$B֤���]��ɘ ��ot���ݱ������@DWe;�%Û.�FqN���Hݖ�[�~S�M��L?贁bEK%��&?rNX�Մ��!O�v���hVau5M���ݝ��!x��ݝ��CNp� �>�!www9��癹�c��j�wuws�^�t <d��
?��e�w�UӃ;�*��7r��ا�?��LA��ݕY�+ς�!�ʝt@�-]S��7=?�T��~KԺGV�%�omrt��j1Ͱh�!NN��v�6��&D�tp��{��Ѩ� �%��D�g��\�ί�*i�ַ�`�=�����r�:�9���?��LX+��QWh}?�����om�A��4��D����  D<H�sڇ����	�B�,�/������V���ABsZ]-�/�m���@��vlB��aG!I��>���ݖ��G�-�u3"[��	6�x�q���l���^�o��@��.��P@])qO��3����ZD���.����3�Y�i(�`��@;���=m�5����h�ݟ��OJ4�'�7�*��r?9�ډ�_�F��閪<~d!����d��Oj�\kJ���������fJ;���"H�"lu�>�i4��B_���#m���ad�6xc�t��;~��­n���8EX>;*�9C(����>���n2c'�N���d���\
��#���eorR�B�WW_v.X���u����'�����r��+!���첸ؗ��5W�9�zeMx��';� ~�y_m�Z�whn�ğ���ۑBj��@�K�f��M���P�%:W1��+ט��9ײ��h�� B����	� ���[��Y�|�c�V\�e�!L&�h���W7r�D�gO�����߄~^_]��T��V��I�k�W���	?ZV|w���}*
��d�jR�xG����u(�;e۹䇎t���B�.2CR   �ᨑ�WQI|����&� ;���g�2��e�[�F��F�V�YE�8�.�z�Ym��m�Dz�C���P��k~�y�e�:Bk3"��a1*d<I��v3&�)�w[���S��g1��q��V��z�q+ڶ'��Z�(U�m�rm��/�1叁�{�C��'1�ΔH��~5}��>��,��g�|����b�kV|=����ʚ%�t8�����;{%�i�#�a)�����Z�`��B��e�Y@@"^��*F�切Tbͦ#_�w��u�NC��t�0V̓5��G�2�4LL�F���o��4i'�1M����x��}�c�~���mۯ�Ν����1
n�J�L;`�_�~�Ǡ"H�����A�Z�d �&�-�q��k��Q�>6ѯ�y�SyҰ��r������	U�j1�4��{��a��4N<�Qm��&����g���/���>�6H��P�2d����s��n�riWc�Bj���F�$�?���/��5Ql1aϵ��V0^�����t"o���d�|g.�bI"��,����T0�z"��Q{�� y9Ǹ� �!��6�E�(�$ߖt��k�+�A�Y�#q��rd�
pAV��N�eN�X�"�c��"��o� �Y�ٖ�R�C�&t{=��3�AB6�E�N��z�Hё�����%��;����e߱������ݳU�fb8t��`�@�8���f~R&��]+ĮK����\dp0��_�i^6��i9�����q���_w�H�j��S�V���f��<rڜ�����N�c��!e}�N�j�;<����F��[8j i�yI���\����*Wn���I��C�n�V����B|Z,ڬ8��v~#i����k�W^�9�~尨>���	��\1)7�ﻟ)!�}�g��sN/������oĖ�}o�!��G���o#��@v�ϥ[�໰�qۮ�����P�#T��]�gR������^��4(Z�%����P�#���U�M6�Ƹ�]�������#H�=�pb�:�{�z �w�7@���H��hF'	9ZuX&��C?��D�,�,�^�mØ�d�@��,Wcl�;$��\�m���.�h	.�H�	������OU��?M -&=��m4Н.�KlE����lLd9�I)Φ&BpD��ɥۥ��k�����L�s.��vc�b�2�^x�����oXK�gn�Am�f�&Bs�-�w��8
9N�<#պ[��/�G:�;z�r_���""��
�]F�˷����-���=�m���c�+��p�;
���ڈl�Ғ1R ��W�	HG�k��da	�� �:��~UQ���Ǚc�/z���T�H+E��/��;��^�m��
�E��y(�}��#�Ѩ1P�2� �z��� �Q�X����x�:5�B��ri��HLv���!���J@��e���� "oɄU>���|Ϫ���іF���pD{DN}���֬�$��קq�N�������>��%�5�
�(3c���kp�y"�C�w�M�SR�1o����D��^O���0��������d�$�g��3��a"�v�����^u��:�x�K��0o�E%m���2Ҁ�fOߛ?��3��џ�d�m�I>c:2z�hnI�ǅK}fְ��S�F�qEeo��w�WB!�H��.x�'�{�nC-7;��>m�skD`�dZ��
Lޤ1��a��?�<_��O]�@���X|-�ӥ�{D���o͡Va�\�t�3W�.D?L=ύ�[al�W��~ֱP��C���\�������\pU/L?���=KY7�OBن��HH-�D��O�F�nE�����VLLo��aUT�h�Y��+�fv/���ؗ�f�Q|����o��\²8�<1��S�W|�M5����hf?�
���� P�9��1�$�R��4�@@���7�P/{���	�8ת+���(���~������}s�����R8k4}��f��D'j�A�N�*��Pj��ط5��W,��bRb�&� ��LT��Iz�n	K��?>���X�:[\\ K���ͬ����}�`��,��t����N�+�$��"����(5�i����;�8ɒ|�h��[1�ߔ�F���
�G:�EQq��忊��bX�lx
b��sV����D�����Ez��^�,]c�T%eޭ,�j��/�8���4nّ�]Q��$������ċ`�]Ԅ%{����kG�48pz�5�J��GX�y�dɲ.�'�I�V�G��u�mTS� �ЕU���(����TV~{�dfm��묇��C4!_����&hY�ԇ��D�<�Zs��f���*�C�}�����O�/�S\��*���?�2�}à��q���Q`�N��~=�-�<_E8)�@��Ȅ<x��Ի��^�{�~�$7��~�HZ7j������p�C=��w�����`��'���'�^x��$g}f��UI6>TN���ԖyE��?�bG�@�*�sQ�;>Wc��X���6����ÛP�!6R(=�v��g��sVhx��`������K�I6�}�;㻹��;�_�7�r��*�wbg����X�<w�[�7;ǈ��;��/��'�}o��/�\�� ���~��I�kg$Z�͐�4�9�%"<)�U52<$��NR������	��dM2�� ����0�t�3{����x�c}�&��-c4,�rr4������u1�@
#HH\�E�H)Le5ܣ_vc)
y�`�U�����#E��]y	͇#��)�\��$8�PH~"5ħ��τ����h�������S�N[P���eii.�;���R���LL����P0]�(P�V��p�A�tn٣�7�p�s��RY�qv�Ҷͽ&	�8
�ތOeH]���賑�.њ��y��oO�*yZ�.ZK9�L�IX��gmk�5��%@X�A4��C9F�R���u�������LV-9s�g����X��󒀲H��ƺ�Q�\���m�Z��]�0�����2E��|�,,÷��DX�kt���Y��q��H������i,�|�|��x��O��LQx�'��i�>S
��i���y譿1��ñ����w��?ɬ����$`.t�z��v��N��wx�����4~Kc)��ڈ*�|�3���w���On��[�%璮.�C*� ~�\�`�M��X������W��<���|Λٟb�"G�Q�>Iw��'����2n�$K9�p��H�^'NC�ޕ�ꭻG�0߯�������^��:v_f;�5+���&ʖs]��7�^��Ψ�,���b�O0��_b���ͧ�s^Ɗ�4
�?�����c��[�WZ����1���uZ����^Bg|J-L�~S׮�P�"�ѱ�$"Mҫ5��8Ȅ{�O�FQ��"�< �p����CJ�Vu͡��%�_�\Z�A�śt?��g�X�W��GM���v;��m��h`���g%���,�6t�I�
7��Z��5��� ���1[�9�X�F�껗R�*%+��d�߫�z�]�{o���y �h�̞8�\������	�@�OW���CX���6o�0OotDu�4��Z�r'��.)?>�]�����ƪg~�	z���c��H�C����Z%pVO)�-wh(��6<=�L^�+T�QC.cd���X{��A,�.�6g�R0����T�u���@Q]UULs���W�U�#o�s�p���C��@ZH�T����c��ٮ�1@�v���|�+����,6�!�<��z0)+�l6��zS��]�q=@�� �Y9ZonA#Y��r����-%Ltʯ�$u�]q���;��y�����ï�FM�Bt�nO����4�-�e�6'7�R�Y����
��O�^�s�
$B����°3"�7a��]~����,�R2|L��(I��:v��p���d��U���
�gz���^:��S͆�ď��b�/@�AgI7Y��a�}3��7��l7�ܾ�>Mw�7�&��ʂ�Or��w9� {V���[�y��k��'R��; 0u3�b����� r�\3����\EG��_��.8�ǃ=���c��Da�3u�����)����З�D^I��a�n�d_��ӭ�_^H�>vc�(E֗�d���NL�`�~�;粁�#E���ғ��r�Ԁ܆g%�:EE��-�������S�>�����`A>�������(F�^��ࢦ�X�~��5�>Q�/�R����"�1��!�}��l����2�|��>�E���$�)^�/gt�C=<"~thS�B�r�`jaV	+�v�S����4仒f�?\�Js���;AhM�wm�f}O��O
�=DP�>��X*���m�p�H��S�l�wލ~�ȓ�+����<���5_�I)��]����,ʰ&��޵o�7�l�6����^��Z9BÆ;��ec�	 �[^VlB���W=o칳�j��T$oϿ�3�qC�h�~��F�^_P����1g�b�=�P�{h��h�v!��vd��2*d��m�o䰱fx�%�ސR��Vnv������I�w�4!���<S��IM��_�u��˒5��O�]���H-rj8�jJ M��T���Tl�eW�=�����o���c�?���7(+VrT`=)�u]za�֚N|��M`�m�)�)4�橖����2`d�ys�̕}�h/'��4;�x+'�U(�1x��˹�'�J�+
�yh�"<>�gϹ�穻��Ǭ��íwiD���g]�a!�p����l�(!�ԗ,�Q�+�R��\ժ=%[�UF����v@����r�ڱ����H�&�,o-J�V3?.k3�q _?x6w�h���E�NB��7�����|0짨����5T�Մ>�u4���رr�V�m�t�pkO�7B�A$r����dh��3�	l��+����8���t�M+������P��(!8,�T�#�?S2i+�]R��ȸQ�g�Vӊf#K"Au�G%�p<MO��N6�U�����.����aeP��Kŉ�/{�,7��߱�03�$cd7n1����U�"�U��ǚ�z}��ś<��FL(�h�:�f�|�Q�ܢj"��D�ǜI��@�^�X�u�2vN���n�mYT�X`��U/�����޶��`Z��#�{��b��bq��I�Uy\���sg���k4nq9���S�eC�P�$�9�z-Y��B�s��DO��������0�;��g������ļx�B�I�'�d�[8�/V��3#m��$�zS�Y�n֡���t��[�INM'�)0�gx��;A�H���к�ϙ��<�T|9��3�*o���WVX��B��M������[��`ϸ-��"�p�e�M ��q��_
Q#�7��I!����|�L6
>�bYl��G�o���'��L�N�����Ŷ�J´Ugm'����������Z��; q��ʌ��\ɪ��\�pR/ϥ���D�!67?/���pv��}Ŝ�OQ�����|�^%ȵ���>ȋ*R����#�cx��b��.�]��g@x1=�3~�(��gr/�c�՚����hí{�V	RT�Y���銂,C�zn�U�5��G�E$J�Ǹ�-ȯO�GE�$����#]����D'Sp'{?i���=N>�ƐI��+Z�u����#�[�R�A�d�WJ���ؖa�;.	sO�3�G�U۹��f���:�j��D�f�'*��2�qpԈ�3&�a�5���Pȃ�x��30fZA�vA��&ΌS'�	�}F�s�Dd�Ц�R߾�&*��B!دg_:�4�����7;���֣�&T0uZ� _���me��Ч�>���_-���7��~bN�i�^_��d�T�A��g��n�V���bP�'-+۟o�/z�h�,�)��*k��x�Am�����)��!��,I�=9�D^�۳>���rM6ڧC��1l?�$k@�!�`\Tf0ML�*J�x�"ʑ F���m#G�4��G �9I��J�Y�y�m�rN�㍐g�;Z
9��}jf��&�1�ƛ�u�g�?�V��bW��)A���3!՞�z�k�`�i�yM͊!���o)� O��p����� 	1a�V#�7�qJ �<~��jp�'-�j&WM�}
I�P����ZN; ,6O1, [�ѵǐ���o�@�$��?=1''�"�l��S�\YVw����?-����fPXjC�z�mfh�Y�[�q��
ԘqR:���5�H�P�@g�w,i_v\L;�f�N��|�UQ�x�;�s�� �"Hݟ-�c�HR\0�[2�T�� ��0���!,bb��^�T,u��/E����^��'D���%�AF]��2Z�2��T�|x� ���KP[�4�Of|C�����b*�{�����"�[qo���ض���M��I��y��L��S8[T������Vh3C���s�H�:O�g��:h�=ʞ� �n�,���Y���`DTn�M2y��[wGH��r-5�.M��o�o�ǆ�!�fSRAԣ�w�ixx�]�g�н1�Mah��QN(�yVi}@��-G�%��ۖt�͕tQ]̡٫���g��zvy��XI��K"���L��7�
 ��S�bD]��CL���Z�H"�����x�Y;��Ap�:�͋2F|�� ��%a��1LN4��CF��}(������*:�j��J&A��=k������[� ���f�z�Z��$/2�9,�}/�f�x�t����[�gV���}�#v�EAb �n���":�0�i�� ��[K.���l�������$�7y!��p��^�YOv;���eD�2~���zu�,`�Bk����$�<�r�7?�0{������У�cє��,��z�sӘ��E�R�܈��%�G��X�ƌC�";
qw	����x���ۛ��Z. &����H*X�)ai�Q|���[����_
È0.�v�7�n���R�������Kזּ�%�
e(jM2:��E����j��
%N-�Ch����i��9)�we��}��hevGE�Z�&���Շ{A���0���ׁ0�_M�La}�<�
c��(�}��I'2>��x��~�`�� �8rx~%��7�*d�t[�dơ�m���P�3c$
s��_ձ{�L&Mʳ����}[�΃)��<	�%mk�cc���JB*e�xGr��QWE��lD��P��y�;���S�uͣt��P~�g�O�dF"�Ŷ��cz���|�f�;0�����7�^�����_II{R' ��w���~{x%��R��6{��Ԏ�}��80vwL	^�Htuu�d������d�9�>6��~zY�����ϿQ������}�nV��B����|��GhΒ�^����, 2�S^axL��J"���{�=^}�;ܵ�^�%נWD��e������3�F�އ^��6;=:���KZ/�VB��
�	�Ahk5��k�`��ĵ�n�� F2b40R]��~�A���XA���2PV`��&(�+
Lv��die�����K(_۵|'�]�i��<+
���*r�0�n�p�$G�����gLCw��rRG�,ꦕ�T8̬��"t�Bo��	T�M�a^�چ�O�Xp�m���"K��K���d�Nd��B�8�n�K��n�^Z�Ѡ�0�� �X��ʲ��qB���1�͸F�B`%5ddX(�!y�	�ݱ1���M���)�J�̱R�$�L`c^|�a��␣�}�{���+��d��2�������U|9����-+@:����bjx�յ�!�l�V��Z��k�>��3���5ܺs��Lަ ���K-MUoh�Y`6$Q�D�� �_|
M�r�(9��?���Ҭ�b�f��a� B!��brB�-8Q~p�5c
3K��'H)c�a���-ީ�u���Ɯ�P�W��y����;
g��;�/n��"�*k�њ�������8^
��^��>��6�b��N�w�4*W=?�l�n���63�4W�e�z�;Z������%]�㦣�3�Z�����I��Tt\m�a�m�dz�.l�~f����i�7��1M��k;
��θ7ڝ�<�{��ӗ��̸݇7�ö���Q�����@Dwݏ$�7��� ���F�GJ)�(�AG`L��镡�s��P&��W[�I�W�4��Gq?��u�N�M<��$��[-A�p)F�%��I/�<H�c�t~�����Z�\�!G��P��]͠b��I��3�\?N��>�Z��G1c�"?싚j�����
ʄ0�.���k���VRM��P���S��r���!~�d,!�ʰO�'��ʔR���J�1����A��t�h���i��Tv+��*�������n�3��6�w'x�1ڟ�i!4��i1lXѨU���S��V_�o��Z�b˘� lm4S�K���S�|�{n�b�eҘ'J=-o|���:(*�8�����䀻lt��FU���B��b����X�z�]�O��x5,�P^��)���Ѳ��|�p�^���Ak��̊�
x��C� �yD0�T�V��28fJ��-NǥP��'J��B�c��lk����J���D�2�,�����-�跋ׯ�O���7�܂�b���m�hJ�_6�C����j[`,e�u3\�-�)��eNEDː��Q�q�����t�dM��lr"���ND�7��:�z-�A�^
F8t��R�2��1�T��M7	n+3���
� ��7^��g�HH�� �+LM~hwV,]6�K't��-U�E��
�I�O��Xl׃�Ĝ�tg�tm�rә&q�!�[�ҥ�ĪG
��)[�������ͱZT~0���N�SօTTL;���B�-YF�r�ɓNE=]Jrf��v��?ST���kV,���$$���I,_�	�2��y$�Jͱ�G�c���I�����?�ǀ������B��4��N�����9'�J�Z�
CK���"Fk�E\�l�|i���:�1�W��g�_8K��[��\�� /�ˊ�&��Nj/E	yhv��C�Co����i�L�;�g��.)T���O��@3Ǫ� ��JM'\�$~<]���LB�lK�r��6�VPٗ[�a�h'?�Z]c��N'?!�<�����Y~��*o����[>�|`�1�I�F��.��/��VLؕ9�@��lw�K�Û�k��[�G�<�uǞ�@۱�,8����N}���)�)	H������* t]��]�(:���C�5�6��0\d!If`9��CXr8��E8N��4�^�2;s�1-��w��O�P�c�{���aF�d[��tR{�deU��z@� JѨ�K�E����C���ڿ���Cq(m�����}�7�Ͽmp;b������J;ǍY�.�����z�������1ת��4��o�sfc�!4B�#�d��w^Lf��4�Fߕ��~\��~��ފ�xzccK��n!��������r�aJ5 {�k�?���LSltdu+3|'�����5��*SP�v>����w��8�y���\93	k��.] �`��P����d��~���O�������%\���^�N�$�X�A���_&��	>T5��q�X�)<w���"&e�ђgl����sG�}���=p�?T\����1�c��� {����p��y���m+�,���=�Qح��j�j2_ϩK@�v��w>���ުJ��!���]0���bol�F$H���3�������^�h$�?���J�j*�K��O¥XnH�t�s��ހZ�����F�3�a��b�~U6~������u����6F��f��=�[K����ӟ?�rzC�� a҆�)3&���m��iW��jD�n'W9��[��	��뫙�����3��������i=a;�fK�q�ځ���ǅ�����D�i�˯f��������H�Q��:Q�pU�Viz���W\����8g�(��_V�q�]p�^�O�1�u��;t�_�',��e$��D¦]=L�Yr(�݅5qr�4Z��5�t|����&��M��%F�� #�٠��Ls���TY�~j̖�#̫��~�P�	���"�S'+h�i�`��ɝT!c�cj�w<�[�e;�V��Ѩ�6���i:5X7�Ɲ��5Q�^Fo4[�ƣ;�j�ǜ��y��-t>t)g���RZ�����5����hr��]����֜��s=$�c����c�N���*�����4�T����i�ҿ� _�U�v0����s�y��t`Go�^�"��,^�R䋪�J�D~�5Z��cJ�O�s���Fs�t}���<S�q6j�PU��ZvϣC�"���fL-\یx�Ji���~v <��{SB��m��,�L�z�]���#8�ӍZxSG��\����;8�� ��C�.
#c�%r!�$��l��i65�;2mP좂I������TkR�6����A=>�\�@��9���d�{Ze��ܚ���Q�����^�`�(TS4�Mߗ���5���72.�ё��^x74ᥗ[L[Ģ�����wģ*��qg@9k~��:���8�/n.7��3�T���� J<��^�r ��Eg계oT�F������B���J��UT��������S��b��ێ�x]��jj�������%8W�S���p�j�|��d�l	\��K��a�/݁�G��SZ:��B.�P3�2���7uK(+�l9���Y��Na� φ��.�w�>���ZBJ�!��CMhchۘ>�0y6~�X?�GȜ��)��]X/n��<�,ǫ�Q����q���f���'�p6���a�eX~_��t�!})79w���S�
��χ��(���MV.�;&c�<�k�9�й�r��T�)�d����f�|��(Z�|�{���ӪϜ (hr�/Z[W$)���ͿwVu�jD;y�:�
ċ���J�z^At��fSdW�8�N�=��,Ssb�����8ī����Kv�<!]X��D(�B���x�q�Y�� U����a:��4@��Cc��Nl^@������5qq�/6�K����F $Uz=�e��S[���|u&>2Iz��B���6Md�����p�j�n�*o��4Vl\d�x�7���ע���Uc�0��&���&I�/zM���g��z:�b�������%��^vF��Ԏ�����LԎ�uF�a�&g��~�ù��uޅ�f�uP}(Ub_�����t�&���a��#eN���*" ���a�'XȠ'd�-��}�IL�D$��h��'?0Ɇ^�<�^;ZД(~�S�ݩ���r�1v�,oA�[��e,���h�\���%3��2�I�9��~�dع8���I�D�^��G��<��縉1�b�C�a;��z�Y�ˣ�WW,�ћDW]�сl�W՗2�D�$��r��x(A��Z�w�:b�8�(^� ��_�.�a��i��0�n�e	�����8� ���P_���Bf:a'+-b|y�YfeX_�2¹l��"#�� A��տSG���j�~'����#��g��!&�_v�8O\%���͸��ݑ ���K�}=��Cʿ&�#6h���`Yܜ���B[M@Ք����c>��p�3^q_@jv��p<�ס�ɷn�4o��X�DV�g�^�j�w��������׸#�_R��eUCW������c�^�oE��ڣ&��y�&ű�я� V��:�-��� L=�;6�GZN���y	���F6�%��T�-C
��b��e��^�4f�@�|�$����-��������ΰ�;�%}ؠ[�}S�,7t�ov#|%Q��	��_�7I.Qx�4aD�u6�+����xnQ�h���?���\��"�&T,<#��EIq,�OD�0' m� )�n�<���K�.����7c��e���q6+�N��ҵ����d,pƽ��PÅ��B܈�!g���6Z�Fb�K�L"���
6k��[uN��E#D���*)��7��;��3ft#�a^S������<�GH�3�.��B�@�-�|����%k}�O�x}���ӓ8��=����z��?�TZ�D�I�������X�f�3괨P�|�Ȱ~q[�^�!�A0�)~{�`��K�}����$��'\�B����wC��
0*o�5���j$�Fh]0��D�.M>�U�{_����IÐ%���7Ʉ��}O���!���:w}��9Op�/�0�/^Ɠ:)�8�g�GoQ��}EO���H�����9�M��u ���O��m ��]��0�^B�g}�m���=n�-�(��ݦ8��L]_�,u�a�9��r�ϖ�7�Z?���L��<r�ѓX����ª�|���0q�APNd,[q�wo`G�i��2D�� >�� x��9r[�dǥخ�3M��P���t=,�~7@H�^,���^9�@t����PawT��`�د�kϋ�Ncz./��V�����Q�Ϡ��4�5�og�㉑�����p�����.YƯ�L=]�va(
���Pa��AuwW}l7B���OL��ߒ�*��| '��"+=5K'.��4�v�U�-D#�k����=7p]�x�?O!����#�����r�-�u�/ڴ"::?A�]��M�b%.:�0��>]Q0=���0�G���~@�pТl�=��H}�����upƭ��
�Ѓ&��f����|X�O�!I-������0�o� �c}�*��-d4�H��X�ձW�ؿ�֢�H$��|�����Nn��w��d�a&q������NK�
���t%�������ߝ�W��^.�&���p���rM:[��B�~6�{�w�5,#�SO54�z:@��g)�X�;����bm�	C6���i+ĕ'�5���\Q��{n=�O�1�T��9�N�(�Fۈ>M<D��R�7}nT\j��z�ҌO���.�PO�5�z��2,)@�(8� Y�A��}�o^��9�c ~���$���G�.��l�=�}�	n�D���Y�@I���_���S����〷F�lo�	�$�Qx��C�"0��4�
��V����c$7ɸ4�.�$5��Px� x�V,Un�\�a�&�{SГB�d[~і��J�uG��R�_�wx�>�z� m�[ClzY�j�7;���	]!�,_ˠ��A]|���f	��Ð�BGjZ�n�������R 0�����NYvO��ɜJ
�W��k�;7�/���MK+�X���[?��5)�l��9ިl�+#��.��@�꺤�2���q��N��W��4.28h�VB)�.̅����޻a#�^�k�Q�����_Oo}���"��&�͚?V϶`^� M�bS�E�S����v c�����ܳ�~1pG�z0I�sA���b��ל܎h�Q�s�ޞ�k�Zku2�o�T�kɩ����X:�\/�,{��n=�,j���?���A�w͈���S�%�gt*9]{?�t%b�nIgc�,�h�k�,���Qp���q�$��@�ɗp;��c%����S�ԯ���e�&�d'"_S���N��	#4_*���L7q ���F,�D������}���4��(��d[+6�UgМ�-.�	��T���I����ז)�t ;��<#�.M��Kz���{X�9�:ׅ��US���"���u����vP�fi��f�lɜR�,�}��]��d꺟�w|4�.ԅDc'�L��@m�,��&]����^���|�i�c�R?���$��i�>fW��=T��K�'�S����|�0�#�vx1Y<R�ݦ��m��<�8�d8�&~W�ިA�]�e�,�$��.�^H�xd�φH�	T����)�Gܐ�_�{��ܶ�^9UWT�f��݉#�Пv5w߉��`��9���@e�Z�8n��=��o�ٔ�~w\�Ҹ{w��Ƨ1J����Ѕ���Zӧz_^F���rV�b���/���kN�v�1=��"P�'%��	��VR��m��)a�)Km��¡��������G1�ޮ����VC���0]�XA`I���Q��=5�9B���0���-o��)��Ш��7E�3��nȱ0}c���r�);Ų\F�Q�m��x��~��_.Ɣ�FV�((,��n3T�R�!;:�����xI|���16R��f?6|I"��E�qG!~���ε�uN|�����)��5g,Rsy/���u	j�JZ�f����<���]Vn�� �d���Ͻn��mTE��aFF��O����dH�F*c��W����u���Ilɱ!ᦣ����s�\���?<L,���Tx��5�ހ���n� 6M�۵f��?�V�@j���MW%M������t"���p'��B�#�C�G��B{�R�l�m
,h[�d3���A�y}�Ӄ>��E��l�[m�����xE�������9"4{N ���Gh����_���)�KbMPEP�@�2�)8m�U�=��7��zk��K�B��N�?~ݔ0~��d�Y�U�(]^��o����*q�ե�s�b�N��.���?����b��d�,������&RAW��� ���U�妖da��3d�u��Z�!�C	l��U^��|�C���:�7r����E7u�->U�×��_mk`�(��/.���6(������u
�J"����a���:޵$�M���k���;�Ξ�f��gmݴ�TPݎ�!8.E\� ~f��-��=4!-ym�"$iF9�s0A+��5��Aa��ԍ.��V�`�3Y�4�4K�J-<��O�����{��	���o�F�}?�21m�]@�t����+��7Wwr;l������\���(��H��g�L��a@�Z:���ZgX���d66R-�s)�M��u>��ld��z9�����Q�U�`<���:xU%=��DM�ۭB��U�.|��C��y�"{4�ۨ���W��?{�d�J%��(�<�4����$J��!Q]{���U�(�K�;�7�=&w~�X��&"9ӊ5���Or�2�*�h�:gי�՘F��y�끅��v@��o��\Dc�VN;��ӫV�L�7.�+ы���>;�Y;)e�Ɗ��`-u�{����r;��=2�'�J�B��D:m�J����4Htki�,�0^"3��t�U��b��Ӹ�Ջ��`�k�s���ى�PPA�aJ�Wz�!S��E�J,n�μ���b,�������w����V���d��C;�)dޥ�|z7M2��ͬz���-�t9lV׷��q�QŮ'�o�is�N�I����rҷK���r���o[vļVnF�X���G�5�)���c���&���^�M5e|)ӦO��Jѳڊͬ���M��r�q���[�-_����ΰ ����b��w�T��X{��C�k	{��<
&�,*�~v�4��᢮��
u=6�כg����cs�d�<��ʞ7'V5UGC�xj����mcm�������v]S�|nk�bٔ]ZO��+^>�����?u5���m��4�q�j'��b�y���Zb�2/T«vTo�)�v����#��EZܼ��1�c�����|p�����V.'��,��l;R�2��M�c3�h�q�K!�]o�v���c�Y,؂�#�M���;���q�)��(Ex?�ִo<B���S�=P3J'��4�U���!
�}ղ�k!#�Y����]Ms?��J��.���`���7�u�r�HW�ӻ��)����j���E{��S�>)"w�$컙K�� �	�Pơ�Ϛﴴ�e��+*y �4V�k2*&`��\��̒�3m��a��_9�3�C���6{�hV�F|��`�H�x*��?�(��J�J���Ɍ���8qp4d��wv��#B��;��vl��z�z�޽>���n7�ι���|���~^ו"��.�e���xuG����.H�z�^F-Dmh�䰬�f��3)���=4�%�ܣw$d�s���s]p��Vs��NZ�ה^zD�.Њ%No{H��v=�]B+#�|�o��{��~Yfk�g�X�/x+���$�\�W�������]� ��{%-�;����Rt+v� Rze�����N���o%�[���x�K_�Q^B|�3���;曳n'�I�BA��U��/�O����� *�>����a:��#"�n���Y<NI�y�%/uҰ����{X����N̼LU���r�>w*c<����i���7��U�t?�.��ߡ�<�y�&D� ��8�y�qg`G�r�بMЮ\n���E\��
؅��)���wt.(���dZns �_��R�cEӃ���<=��}�5��p[h��|�>*�qg`�҉(E2wH����o3kXM�U�-�X�N�Ƨ[��+H~�����ꜧmj�:@�ޓN��(�>V`-N��q��������|�1x|�
 ��1xz�W�+W}��|�8���:x�VтA�rEu�U�^�6O�99��i/YeEs�SUG�e�[�!6�9�/��I�TPyK�v���52_�O�ȧ��ܣ�P��:�M���~}��hGel��'U�@��' ��9�� � wt�&��[�Fj��
{�߉o7�ND��|G����v፮FMF���Stը�ֻ��$W4D��MX�?�%<����Ca����\*�,���'�	3e�7��
q�f�*g� 
�4�QL*���[���?W��<��`'���Eͺu:U٦ni�;�i�_��$���h�鸙���L�Jw�dc��2�����M�v�|�|$5���s�2x�9� K�LQ�����E|��Um�{:_6ld��t��72��m;'p���X�"�n/��ǉ4<8z��d��\�>�j�RSli�x����T5����!D�j��q;�#V�v����!,D�X�q�ǋ灖A^O�y�e�JJ!t�r�7��˒���&Ȋw�����_��?�^�U�vh��I�HX7K��L_@+�$�����\�'Y�������-ZS�����AȠ�^���h�ǑK�(�o�wenX�7�V��A�����0�v�����W=���W�:�-9�3��'��Zzmn�JH�d�8MW�{M�o������EP|��œu�0@�9��8Z7��8����9�_���}��v��ֻ�z��k�{���p����KY�u6@����v�V||~��"��Q�+�͹o�<=� ��SaC[��^	�Ox�,'><����x��^��1s��]� X�������r$�c��i�F��.~��Z�#Jt�'! ��r&}Mc$��W������2�jѻ�ז2�P�w��/w�:�U�Q̵�hU�qK$RS����ǼP=z^�(S�k�Q��v��J��d$;�Z>�{�ׅ0�R�����2;@+����(	e�6\ry�:�|�|��K��ś9�pO�WkP_�+� ׸��B�:z�A�{!�m�m��vn����"�]o�h�eD�G^����+w4�*�䶽�b;6�.TM����d�?��y�'��WT��Z�&�'=�Tr��[S_�����FV'���e��00���(|�{Ba�χ�$�;$��G�jYD����vo���)Q���ː�bN�sl����j��2qw���I�d��g M2-�k摵�l>��F��K9����6�tۋ��IJJ�'�w����o��+_j4��,�E'��߼O_�!��*�C���4��B?v���7O���:K���=��U}k���c$˜YA��-筀N�s�{���u
,M��]�EDPc}��<�f�J�I���_��8�}��P3�T�?�/��43E߉�!{ɵ�E<R�>�TkVt|ȟZ�%��q�םsm\�j�t����^7���`�j5�	h>f�5�6�dI8��s)v�
��@)�����iy�3"ſ��n+Y�k@�K�]�Ia'o�DHDUb��&S�
��<6c��������*^Iژub'o�-{�U��V��M�Y�T�|)\b)�-�[��U�"p�_,�%�D�eI�߭�=�q��1�qK��F���mQ�+&��m$�H��	��b�J��a�y��t~z�[���wO|:Q�W]��LX D��s��%�]���zz�׼�Rq����5�	䜄���l���vg����5���d[�e�_ȶ4Ǘ�{f}�*B
��tBO�ڈ���S��d����m{I���=:�
�o��+�q2Fd#Za޵�����-!�_ӥL�� ��q�򅡅w���좌�/x�=)N��t1N	��{�A���S����P�o|�T�r~�Z���C�� u&�z�阠��q� 4b[���� x��e#��\b7c>lDw��M�^:o|A5# �YZ=�ա|��	��Ș������T���%�V�lCo�}�[|��0��<898"/�кn��,* ��w��11o!W}���Җ�o����h��,��^�Lm��$��n&��qU�+j���F��Zwޯ�K�d{B��_��7ܿp���_;�K(�P-�y��"���'����_��8�G���uZ�lI�oG��?����(f��1h���gQ?��y���vw���_��%	p���eS���%�_?���z�e@����7�ft}#G��¦/o��'s`�6�����n��f�2����e����+7���\?��D�߭�|��ق�_N���1~;b��=��_[�h���s�q}����ֿ�#V0��X܆��m�}�����I^�'����K���������|�c�h��K�=��{&�gL���������{3�V���|hi{`���x��K������Nk��l�������w{AZ@F|��A9  <�~!�ۈޤ�V��q)��ف�ՌQ��B@%o(c
`^�봆��F����PR9������#��w���-�O
�k����=t�	Ӥ\k#P��7?����Z�0�������+}ӯ'!��B87t��.pU� � �d�>j�~;|7_-�. ��2����{���Կ �ҏ��g�ڧ�ŘB� ?S��6�,{2�֮Ȁ�����7V::{���N�����Z%�b�~���,@�~_��|�5�.i�x��6���b�m3]���u�-��缛��e8����A�+J��K#m��ߞ����~3�����yu�6W��AW��i�~>���OTw��7z���l��'T����QĻ�T�1̛o��	��`���GSenHJ�w.{�w�E>�k&�䢹�.ݧ,����o`>�� ?�@�?�w����zP	����>�s���Lf�ض�+�5�2�ik�j�9���jqF��7�ʧ/d�_np(������:+8�ڢD�Q8_H`P���펻��`6�p�
��5�tthS&�3/��_����3uaм�<cPI�]��-d��������O�ߋsi���	D ܃%���\��/�DZ��;��;p�Bn���v���M-Sg��o���T�]��I^؋�m"��/)Z��$��gJ�A���or08�;L7<1|0vW�k0��k8��O51�<�iGZH�B�R���ox݋�!���	⑂�S��S�[��9�ty�]�g|�/"�{n!f��Ɉ�x	9��bP���F<�Z����bO�&��^$�
Y	܍4_uou�櫬D0*e��
އ3R��`~ܞU?9�'K��wIb���g�s3���1���Q�i���!����t���F!	���p���̥��̔/�F,<6s�Q*�-��ۏ/�N\��y驼�(}�Ԓ,���<�=��{ 't���ZZ������ݤ+n��nЀ�2���M},�_Y�aMAJS����Ԯ��ő{?,WP�N�~C����e
	z���	�� ��&x�B���]6m>)�˫���ĪE����"�����8�!�b�
�ڽ{L8�5;N���o�a��U����
��5O���k4@f��^̮��zȒ��5E5C�;�g^dɛd����������Ւ�uN�{����~�W�����1b���ٻ�nN#����!pm!���*�_�6�l�a�yc�������!P�:\p~�:�P���P���q��S����#�]e�������?��%u^��1	�>@0�"i�����]�Vwt�'y��J�ɴ�9N�.�!<�B�=LN|�Ѥ(X7ϧB�D���M�
Q-
	�U�~��]e'�/�u�򘁫�^��I��2�MC� �0�|�2	���́x����nY�C�����Y<f~����R��M|��KX��$G���>q�-[\�}�a�HOɱ��M�����ē��i<�o�7�F|� *���֥�N�f�3Ƌ樂�,���'��sZ�IB�3y��UQc�Y��㒣Bë��>U�K�c�������dw��[h�t�@ ��f��0�������jaH��r'K�A�
��^sc(n=��5���v/D\*�Ke�a�'"B�qWn�}�_$���`rD�+�ʚӨ�����2�������d�M�Nu����?E��V q��s����������2�\�T���FVq� 1�2����������]mf��ù��D��d�E37:`�����g�H�Y"�_��.MXY�U ˊc��u�s5F��w�R�5�ԋ��s��ӏ ��1Q�G(��$���sF$A���<�yhڋ�>taKD���CC�˳��5ouv�X����7��3?ǿ��5���NF�_}�>羍<��CVȓ��끷vu���;4vB����^��h�����t"8ذ*|���uZ�M�"���(��ڛ�ez�d�.�Xqv�s{�󆟸�>;w���0Md��,>��l3Uf�����vU?��T�xA�4�Jw2�5D.K'����C�7+t��!~E1���I�~P�Ȁ�ɴ�Ζ��G8k��~��yg�S�R��5�E��ޣ�=�d)H�Qu?����t�r�p��g7�@/� ��O�G>��S�,m(��:�9f;����)���9
�%t�d"�>���x��;�x<>�^x�H��3�,���Ʉ�{C�TƑ̤��l�R�4���x��J&g1[ޕ��L����d��#'*��
:3�=�N#f6��BN������;S�����R�+��| "[r]�0�s`@�s�'�Z[�m�e`�����O��-IB�uT���r.�ro����������K�ҭ��/���آ�[�����r�~�Hsx*�L�i�<%*�Y �>�^/NJ�p�j���>���+5�t#�C�f��]��DF��1
A~� Ѧ����jT���:mC�a?��P��Fߢ*H	M$���+a��!���A���ĸ
Bh���`�q&D3Ɔqau�3�^n����D�3Cz�R�>�^=�^$=�D�&*�+��!N���(U��e�4�kE��w��)RFV��W���U�pѪݴfB"��m���GF�V��h5��|����mx��к�r��Qv�vmxx�Vz̰�Uֶ���y�@v���6G&D>�L>�nA��ŷ��g�wP�� '�-Gf��Y-��22aJ��r���3�#7Y�wHl�c�n�h�(D�F���dX4KڸMMq�z>�!��"����	ɩ��i�DFῸ�n�~��;ɇ���q�����yγ�*�V�DkԘ�tQɌj	��E%��S�ɻ����V+�Go�{���A?�dP���޽����C7��i2���"��&�k��3m(��*��"��Zfѩo{�i|P���S9�I�3V�	b�+����y�ĖoA̦=y�y}����Ts�a>�xAS�b�����l��{� �q�&�|��|���}Mg][d�h>ř��Vjd���Ǡ5hGZ�O�����x��������ra7�[Z�i���u�h72F�XXI�̕i6�3y����Yu�޸��zW��55�:�
h�<�y���ߪ1�����N���ʜ=�g�U�7�r�wB'�u4���|.��G��͘�J'���ha��޶��4�:�t���f���Z@��G,��-���F�X!b򝟔�#y�
��#>٥����SͩUG{Ҭ��-�[�	:@,�>o+ٴ�"��O���g&��Vz��ڊ��qT�ɠ��:���gT,��~<�+D�:#�9C1wc�,�Ȏ�!G�&�L�	�f�2H4�C#���8GN2�E0�A2`�۰0j��)1���i�Ey�c�]�GNz�v�~v��m_&ѿ��P���$\G1����}��"���(�g�r�_��0�+�eau����b�_;j�r�T�y�'�3�5������S�/�x��v�`d�� �%�RyW�2B��S��5�6{�E9�W�Vv���v>���3d�^
@R>xYg�
���\��!����c3Z}��Rl�L��_�)��j/m>B�����(Ie=��y{�l��sN�b�x+<[���o@?l�Y	���5��%��������	�Z����V�Fw�t�l݋�k[=�eg!3�ώ���;"���E]^=�lJF&R�@1��w���=����;{׳{�k�,<�yQ�ظ�r&�m��=&������`�>����O�D��Q���(b��z�5g��S�'��9<�@xz�U�K2��/�mX�U�dJ���w{F[��L��o��5V1�X��89��ɞVx��^���T�n��R�%0H|\�Aޢ��و~�$���~��I ��\�:.�i�a0��]�i�j�۳/�Y\V�)�{�>���¯R��h?S/����Ƽ�1_�N;
��Rqu��ҽ��Z]���@h�1�0*?6"���hfB�{^�-2ҶbӸ��L��e��Ἴ4�*ˎW���z1A�LM5@�7ܪ��FgZ�8ר8�c��C�����EzM��尞|�'Xq��J�*��}�0����OC=��Z�n�Q�~����h��9���LK�lM��m�w�]�K�6(2����c{���Pa�CDx�^�
�:l�C���$�m#{�����GI.^���L��U� >B@����?n�����pfg��E6�{�G!*�������7j���B��-��J-�����(�;������E�#��^��L����<9y���������Ks�%�Ώ��b���H�������/�Ѐ�z3e�z��/y{x�>�T3��>���kp��@q��K�<.~\%PW�\�o�U����1�= Ls�=mwA@��g�����K35��C����R\��Py���`�$���ԍ������ndR}���92� �~��]�qfr�B*��]�>D4Y&.[wSS�Hir��=�P/�4k�nN��߾ro���id�y3j��/Gݍ�mc.��aF�r�O�1��~�����:~c�b�0p0�Wn�'8�E�MP�����Fe(�wF�/1�����Sو����Q�B[���YJ�@�Qv@���i��PBҎL4u�!v������I�w��L�[_����X�JmH�Z�K����Hz�On�lg�S��,�/YBg��U{-8(i+��q��o��q�<o_c;��k6���E��7ц����ځe�(��3é�-���-Qh����-I@`�*}�-����tP������?\�e��j��o�^�a�h�^ ����x��\_9� 4��N���UރR��]�9�J�U�Ԓi? �l�i�,��_=I�Y�sv'����w�ngg�s�)G�ś�D2?���Cq(˳��H�0(θ2��6@���%���tVt�Vh�8�N!`"��ǹ��>ٕq��Ȣ [(@���g�+�7s��i����$7:�Jt-���pJ#����5u�z���Έ����L/�����0	*2��7RN�Mf�:���9>��;� gܯ��G]t�ۘx�My�L�K,5�G�$�&9��.L)9e�zt ������-R��r�Q(�m�e��n��z|�����S��[Uٖ�j�ϛ��{��A�9���u�-n��H5��S�{_�Xw�&�,!=k	%?φv��ȍZ5Ϋ�{�b��{|����NSm]�f���V���r�nC�}���� ^@1���5HB��o�,�b0��7Խ������_7�dY9���)%����F,(�FL�����|)�7�S��EZ��ZF���$�˂J��$@�H�3��o�Q�9߱�z��,v�`�e'?q�m��V�B��][$���?�:��W�1 .��oN �z."w6�?$�n�w͕��{X�LC��ZI�8)_���w�P�c���6��yN�<'W��CǝG\�[^���� jǝ1�؃�����eA
s�m�(�u7&TU�v�N�M�ꇷ:��w�x�	,�9%��`����L��Vr�kڴ���ns�@{~�:�M���s�pƶ,�����M�SK]{��R�n�A�	{��c�T~�ϐ��_ss�Ip`u���<Ub��K�Wݲ��H&oԠ1��v4.
����{�̆?Mŧ��;+g���۸���"�����VG�$�ҩy��w3�Ͽq������gs��bc�����4�X�3�)�9i�߉M�d���ׂ��B������Df�@�3ᢖR�����r��W,��h�� �`�~krt0�',H�	�e���O��qў�t���hW3@�{�:�D�O��	À���c��?tr�!���l�m�8w](Ff�]�G�6�л����t�0[���v;}w@��bsq���8�v*��D��D�:Q�Wo����'1����Pqq�llj��k�%]ֽ��W���gh;8G������鎖�OA�� ޷M��|�����UW�l3���#�9����87ۯ0�|򪱂\������ꩺ����̛��� �3�n���	KI��cA=.9;b��6P�2Ѩ�/$$�(g��Ǐu�		}4�D%�m�DW_c���Q3�67���Jlw���e��ʩ�F�Z ��t߿��{�y ��P��t�h,���+����/�]���X�L��4�������\��:�
��=���y��j��q�#�1��Spӎ]pv%*���6@�m�؇�Q���Z.�Pg�M��@t�����W'\-P}fh��o����@~��w�%ex�*��]��k�߲��񴇘��Aa ��M���L��;׼J�ث,OVO�d�Jz����Щ��2s�X5�����w���~e?�������}��J�c�Dδ�}��k���)]�#ś�ŋ�۹;�9��cP��Rr�"��N�<w��w�_�f<Ѭ��*P�"���=K����_�b�	�����~�Ə�;��c��z�s�>p�cP�M�V\>%���v�E`����ME��&�������w����������9X:p+ֱ�\���W,;f�'ǝP���p9��|E�(ĕ�oZ7����BU�&�8�&Zw�2�L�DX4D��
�4Re�� s�����d짂JI��t�{On�^Ŕ�����:~K����Ϛ4-�aCBh�82�n��w�o����^2Sckkv(��}48�}L��������-�-����s��SE�["�4}��
�r>?��Y2�m�Y6d'��`���X�c��V�	p��p@�N28�,�m����4D���':���ɓ���)qG h)�ߏc���u�H�nh�ms���+j4>2���B���Z=��G�����iC���6��&H操���M�~��0�v����QL�}ddÍ��T���( 2����"�`d��Շ�(�?�ό �Yb�T-�7-Kq�5`���XO�����e����ޚa!B�y�v��S���S�.b��ӓ�Vk�^�
|?"@ZHdB������s�a)"B
�",�GH��׻�v8�
 b
d,(@��-1��iJ6Tw�c��������G�C��0i)=�	E�l�\o�v��y�Ƶ�����Y�Q!pYD(��2�`K����|d�J8��z-�bU�����¬Q�ɷ�W�v�v5ﬦ�Ua�}���&.�VM�O&nM� �U���Lk�Jo�5�(=t"f/�0��I�mY��P��r����^�y�Xu�d!��s��Xt^�HBpvd�-������^��b�;7��V�
�9�<���w�F\4�2�בF�ʮ`���r������U-��a	A,�u�D��D��U��IRI�����T6�ð�.��Lo���2���Ș�Y����n�jDT-J��4O�{�%�"���j%)����6���ڇ='�����'���t���]�a3dTP�t�$���#\Kee,M�
%d)m�x�Y���m/�L����ccK12�莶�)<.�m�2�����2���2���m��`e�krX�2��3 ��f��y��^���Q�~�<�E%3�̯6���)��gW��T�l�n����~�Y��^d�w�𽾜?0Y�"���qڋ�ʷ�����h��O^cs�X��>�;|q���ՈL����=�Ū����8>.�.�k��yߗ�F��1h|˹�q��<�?�i���0q�z�a'�uL������re;�i�pxL��-)�!���L����Q�i(ǻG�ܲ�+� �^��$U��j7br��>���Zzk��M�Kz�gZ��#��47o����r�V��l��N���aS�?p��ռ"J�@�*nm����* p��N������X�O�&�,t��4�L��w#j �l3[�V#@<���?��9����o�1צOE�@O�G����ܱ��d[ȰldJ���pI�3�����NW������Zݵ[���Ov���˙��w}�����k-Z�L�'�(�� ����Ա%���:6%����,�M��,DN���~>�%*�e�Yz�!�����r��dj��1�dNO�K�W�7���m���� 	 �m��k��!̛W�<k^ �
���냉!+oٰ�n�mmͲJ9�L�:v�8��W��~��|.��R{ٙ�#Mi���1�@�b�A��Yq��#�K�&��8_�L�ì2�P����#����X���ʤ]��B�*^V�l�F5>T����M��=�Z��������;	q18��@����<��S���+\�^�>+C�����b��h����X#���t�[�«���HCF�l�Vn7,��ȇ��nb!����]�X��3����#�%z��Qx��[����yV|�q=���oO[���뙒���䪎��e:�n�1�|o�>�ק.�`m��-"�@|gމ�������fS�|�:]0$T����Ӂ'P=�\�-�����G	��ܘl�JYy�C�f��UE�����tBZ/oHAgZ:�7Ci �; ��gd�|mc~?n��D��z��f�mA�"��I�����~�4P�ss��S
N���T6�#� �6�l���w)�*�vݦ���'�?��l,,��\�#~���g��rṇ�  ��Ey���4�m20�:[�g�u�ݣ�>�w^�N�A�����_��tF�6��%�#*62�6���(���8rw�u��dSZ�������Ie�v�9����7��z����o�W�8��>�;L]am#*�}a��ɹ�4_��U���S���ȁ����Rt����ju~�bbޡ�+�c3�d5U1Mw���n ��>�J�2ࣃk�!�B\�Qf|bگ�򞖕/E�3�Pđ-���|p�f��?+B3K}��V��4&3 -2�� �;���Ԇ�%�,�D+�E���R�����eI�j��VP%5u��Syq�Nث�ޥ��#��x�Q� T�R)��6q �$�����w�ywz�
���s���hBCFR������ ��;�/�g��;O��ɕ��U�9�*W�n��b��h��ڳP�I��=�x4:�u}Ջ]埛�Cn� *�Ӕ��+��0��G7v�U)�c�m�����l�,���/�|��Ѓ$\�CTr���I��=!!j1���-�p ��w��=�lݞsjṵ�\dV#xσ������#)z��-p�gb��P����E͹��n6����r@��ݷ�-X�݌�x��vj,����T�j��ޡ�;��H��i<�)%��蕴��U2R�\\:r�)om�4��ΐ���[XU�n����s#��hfb���R���Y��h)��ioU/���hv������{����Fv4����P���f�,L�I�dx�;�o*�Р�o�/��GP�E#�&�7�V�q��$q�\��;T8]�:���uy�3q�
lݸ�p���qJx���/��EU)sΘВ�8����O'��,��i�k�8��BG Yf?¾���bH��N%OL�'W��>�	+QPM���^cK��3�<�o�_0��aV\���Ǔӈk�Ėo겝x�����g�;)��p�uR-,y#�����]���$w2c*�F�K9���9�%��'{�� 0s�����o*���lUl&��9HPd֖>λ�R�!-�G���sfl�]�_Q�]]�CC4-8콹��xջ�s{ z��2�fggs����i���*�V�Y���Z����X�N�-ci@�n`0��T�	;e�L�̾���O��C��1x1Q�U�;�8�z�75=�g��X���򧜰�6���hnM�JI��k俚�w0K�ҏYW'7�}�ko�Q��[�qgDT��0aQ��� �C�]��8�����1�j�;&	����lu�� bغ����ָ�<��C�W�ŭ��6�ľ�LZ��[
;F60l��ʩ��5�nxF �P�%��#5d/�owR��]
���V$�5���%�J�U<9���ܐ��(�A 0؞DDe��~��2&&ˊ���,,��X�"�*E2��_"r�/��_�=g��q�1�k3�)5��n�y(�~4�pM�u熰y)�vQ��^�9C�Y��.���2Bx1��3xR����m��޳��i�������S��
á��(� �{�� a�}�N�>��SK�*|�,��+ʹ&&�f�@� j��B\����O�]��Eo#L�鯴sng�{]k�N�L�~a��k)c-uz:d3䝄����1���/���}�h?.�Bv����!R��q��5t��ȴ6�w�����!5�ky}�7Ϯ�m�q:����VD~�˕�n���aB�2�w�e���n(��%�w�D�y>ݐ�� �5Ą�)DW
�+K�
��r���J}>ܣWV��(N�/~���#C��8g;_���S�e�u6��t	�錱��P,��G���QR���h��_5N�1u�^V�hS=2�����ҙcYh�/�@���vk��>�B"6��̥!�7�1��ؤ�^0�&���'_�3f�f�e�L�$�4���-��}¤�$����ks`�[��1��aK�^�ڶv�"��ad�M�I�R�%h5�JYJI
��m�&��Z��t�����SSE�j-1\��z��VH��{7JS)��H�z0��XFX��

�KWZ:V�I~���.��$�>|  �k���]��e������t"M5�a������2;p�
�2�]z����X�g����%�BU�㪪��z����Q�ʑ)̜�!jC�a�D�vr�Y%�H�[Jov��F�A=�e���Q8�]+//++�C�n��5'm�-��.5�{�L'V�:�y]`:[�R�dh�$r�Ef�����Ϯn�=�������TO~&��i��!++�ۓێ0���҈�ϑ�c+��[��07n��g�a��g�M4.����g�ǙOSR��h �@�Ғ٤Ծ����o�f���@�ĉ�ONS�th�g��)�B��V|�Bf_����$�ӊj��D|@�FA�LFêު�h`�E�u+X�^GB:E���n�g�3��O����:��CV��z;��=o(���V)�-M�"1Db)bh�����#�
�(�z��94�ޑA�f� )g�����jD2Kx\^��m�T4�Ӟ.���-���w�	H������d^�{2hFW����l�#`��3���,�"�T\��7��fp(7|�WF��<�xEu���"����$�5|�� ��N�k��xK���K��$lؤ٦���]À0d�z�J??xB��o�x)���OJ`�w6U�I��ť���Jn�t�"J��'b��|��`~�6���ʴ(�����������.K��0j�:,��Qۮ䄬z�#��*��섿p��
�F����jL�x��a���� ?�]  ز�"Ȩ�H:�à��:b�R��$��{��M�
F�spZH�Z u��@ԇs�]ػO
�$ ����;؛�stLT�?G��\���c�}�wo`��t4����d�l�M���-!v) <f�f���˦鼛Y�ʘ�ܺ�,����-��C+#��#~!��#��1弫�3�G������-!�����^�<��  �Ur����5?�H��J���h�3rL]�AԳ��}^�KJ4�M��痖��$\���)�������z�D���oqZ�$լ�3�W ���Ko]�������:����
���Y����#����� 1?��� ��hY���B�������^1XY�I_sLL�,��H��x��]##������ܤ�i�-����b���B��ʶ��"_<��3na�
\�
�_�i��k�{}�
�B��lu�NQ�~&�#HLR�i��>�8s����^��M�}�鄙��֞��"C�O7֜���՝5�a�����<��~����o��'��{x��̐]8k|��h��z:�]����ӯ�� ݇�J�������R�٢��n���Y�9��@��/��g8��/%�=R�p�?���#JV��ۀd���}" �*n5��;�=7��r6��O�_�6]��m�p2��Wj��7Ja��x:Ϣ�?�E�[ʇ~�*x!���[�E$�馿h���RU��A"��L���⠨�\�=�O���))l�?X��s��F{�'�������M2��H����3�/�������_���R�i�L�t�~31�Ke�+w������F�n��[��!;�?W�9"�����o�c"5?;�锣~$PA���_X�<�7�e�C]����Ѷ?�|�<�lY[��7���'��H�Ǻ�u�t����_��1]I���"�?�W]�2(�����.1Y�6���Ӫ�d����3U��EF��"3��t�
B���^}�0������0 $�K���8�֣G�d~�ۋ�QUt��s�HN�=@r����xzz�����pz�nS�� �[�^	:Y*�yW�g�z����/��_�Z�S��=�i_!�?)��s��z��N��D�9�_��H��:�����˾{�5����S,e����Ň�]�U�.%G���"YD�K�!�� ����B^2��)׵ʓɳ�(5C���$�)���$��20 ��xF_>DV�~Xg7Ш10��.�c�57p�A:!#�X_�4w��1���&�&�A���้��JR.���'��ہ���4v/�Wb��N�R�5�ͳ��*�]�|��G�^ȟ����Ϝ�����"�Na)4xI����(��m�?��B�3�nSR�����*�{F�ާͥ��팋q����!5�r�J:��t@�1}�ă�g�6ύ�S!{�`�jd�<
��x�A&�w$�(ɯŸN���$����U��X��OΆ}�K���!O��l�(}��p�՞��k)�A v2wTp����T7��d�/YX�(5�RR�Ht�����?�Z���� �*������4���G�?��������ǎ���y�P��W�������Xw��c#����;�u�~؞6�)�/[��\raX�2Ͱ��l��n�c�ڽw�0��Dq7��·�<�9�͵��+`۔*��i�kA�!��ͽ+.����7�Ϲ�;��܅3]��#������/�c��Ջ(%㍳�)a�����N	&��[]���2��+���)��}9�桀L�|ZȖYt?6�Yx��������53���!@��k'�����@Η�� W���é)���YA��Dg��*���7g!�p�,�
6?�;7G������vr0���:���g��P���K��5Y<����n���03��y�/g���æ�t����m�g���oxֶZ�&����%L�w��N���H���jY\�u��U� ^��j
���fQ�o���a�d'n�EH�������l�����ځ������sWA������J�A�.m�G[3Y�@~w�@j��3��OWr��I��Q���ڿO�ֈ����p�N|R�2'�������˕�����>u��7���_\����q\M�?Z�ϝ5m��ʧ���$��3v?z���41���h-�d�6�ͤ�
��5��N~�=���Y�Å
��T����:�|�1s��_m����¼���kᣂ\9�ˊ��Hg��[aJ���]������b�gVA�_����GG�?����;����XHv�3d�٫�k��uqÃ�����>;ׄ��Dg�l�Gw��f][��3�*���㯴Z��8�R�������2~F!���\��U^=�E]�W�{�a\��e�h�� �
�i��\z�<�U!K�ٍt�Y_\g:�gh�ީ�I�g�z�PS��CǧՃ�Ld�Y��&��Y��aȟq�G���)Y���ыbI#��,���sƟ���-�_��O;r~�a�����SݸO�l����|����y�ҢB�}e%��a>�yH�j4���Cd�3-��~/�CyϹ
x+�;��.�0���ǅ�w6��UAQ�s>Gd2XŹ?���P�üx	A2Z�v�3�9�G�͘�L��?�&��f�s� =C��kgP��m�����SO����C�'��s����[,�n���S��g�*��:uqū�%[�AV���/Ÿ���=���=fթ�feY/��7��Z�C-�X�)x�t
ȧ���ʍ�#X#��ӥ�l���D��CT�#�C���nW�>�t��?�>1�z�F��鏚�/�W��K��<$N+�X�Ǚ��D�_5%���~e���Մ3;�l�d���Ogr������,�W�`����<�f��ȟ��3
�?����a���#��>j7,ts���\���{��{�.�*���Ј;���y���qBD��;X�dU	Ե'��;�����)��@�'8>�=h�τ���q{�j��h�@������,�����~R���#�F~�{��x�K��:�W��������{-_>��Ǔ�*���I�_���ԯ-X���C��]JY>�C��g�x �M�����fC�ٟWΝ4WL����>��~.�P����L}W��HP<
=��(�CA�-�.,  �0c�k `�qt�9�Y
����u�_\�3�F��˚�A���库��I�T�?����`,��$�0hf�*(�U���g��	��U~�cl���+6�2:V�e��T�}e��9��T�B���wz�DJpA�t�w��*"�I�zB!���0�o>�bi�{��{����{���IF��1U��<�� ;Q�A'ӝ�Vpʯ��e�`/�/=B_����d��H����r�S��V�O+�U��6xx��6w����au�uY�t�eOJ������8
Ѡ�]�?��D�v��63��b�]'Qs�7��f�qvʩ]���@�@� On�~ �r�������}��߭襠��;	מּ���X|�brx���+�t���kV�$��x�������2�v��B�e}jf�_�]��|������T���P��6�awo ܟ����q]7������2���OxΊ�d[���� /������.@�09�y�	��Ӷ:����3�����ϐ����7��[ܞdM�}Ωt�\��.H���'B]��D������ۏ�
�x;����5�@���h�{������k�ᎉ"���$ZX�W+皱�y�n�N��p]�ۀ �ċ����a����!�xM��)��_Vuka�,���
�)��'����?/�s��P�8����{��mw���o�*�ҝ�D܎��v�l}�|�9���KN����x�	�h��Z'ril�dP{7w��y�
�7�n��4_�o������B�8CO�L�(EϤʵ/SG�/�2ٹ�B�Q3��K�@U]�)�i%�qp��/|�"��I,��X��+*�kA�徛���i�>U,|��˦��������Tz<��=F1oJ��S��^x���vI���`�������ǫ�[ɰ�l��K>V���K�8�t��/S�;�����U7�� ���9�S�����Hk9.^l�G�)�e������83�'�Va�?5��S"z���kg�3D��~h�,�E'4�Q���'DF�RC��j(��\Ŝ��V!{��5f*��!�c�?���,jG�*�����t����	"�F�ؽ���Kdǵ�1�O�F�\IIg<nUxO~g��E�]2���щ��qe�W,+r�h�iF�������ӌ�S�����8'�N}�)+��SO��~��QD��+ħ�G���DD��/J S`}��ڌr�����*��<��`�Eg�������: tu��{��W�܍r�)���udz�p(�uA	�Cg9,,a#>�^�®abvc��pWӿ�����N��Jl={fY? ���O�ʿx�t�v������ԋ?f��cK޹}U�?�T'�zHA?�ӿ�(�X��G�p���9S�f\K�/]�5\�j���~~V��[�F$������6�od�T��p�iE�f<��et�����n�]�TF��d�]�1�W}dA���߅�@A�B�OF��%5tW��YrQ�G"��I�˙�俹����ȿ����MǍj�ܐ�~��_���XlSfJ|��K�c�X�_��Dß�q���/��?��!'�P7���,��G�{TƆ��Z��=���M]n����S3˿�~�
���C��&px��5g�7W�[���>�&w�):j�}����1�Bt?����J��
&��;F�V']�;� <MX����F ��C��¬{��i@�Jz���3�n+���XR���-��E@l�L;vF^[��b~0E4��PQ������=���'z�v4�B���j�a1�Y��G��bv��=�����9r�>����~N��@l�~o�!�O�S�[O'J�0����ѱ�D������=\L7o*:�Y�k;�ښk7����oKY��N�%x��gF �6��8���3��o�k�B��5�M�JǡR�䤕`M���=itٞ���j�j-����u��D�716�ʅdʯ�����g~�6�n��*�bI�=�7"�V�+tD�x����K��ro{�(� �ۄ�LS�����qx2�D�Ҳ�ъ��xK�����VW�����`ZwT��O�������1�\�����%| z���щ�_��;�8�����Vܽ��f����h�q�Ɵgo���3��^���k�.�\9�NO�N���M�DǷ���~�|�g�ʗ]Ynw��29+�:!�A��wA���ڥ{H��h�Q'�H]d;I�?��� ��ǧlnmCF�'�������Ò���j��A�O�Xa3S�|�e~�~���y�u�Y�ț�&� *=>q����"tSF�:VK������m��B�h����$�,� �賠�����f�h����S�}��̨�wG���x�E���wqSg��a0�Ӷ�E�� ����#F��O�%5�Τ����5c�g��q��|j(�t����X�Zƍ v9��Gٔ�br�w�G6:�AV��	%�QB��O����4�I�4���_!{�T�o�&��~����;���=�nv?�[�ҍ��m$���Y�bՋ�W���Z���
X�$����+�q�߿�6��ۛS�l�+�5�^��>[!^?R�o?V(5�4��K�ȕ~8��)�9��|�I��^��s�DIE=<�CT�&��e���$�0�L�ѹ�w�9�k#
!����e���'��j�}��MyЩ+OB�]���M��s+ɉ�N����T���26��K!թ�f�F�`
���g@�0�%A�W|0"�F��D��W�d������Ŷ��uy���`.��~�w�[�g�y�33��Fv2�x�:��,*CA�g���뺬�ς"��L�Ero�2�������˼t ����>y�{���w�^��@�rx\B r�sZ3�Ns4����0�6pW���)�2�	� Z	�	Bc}U�u���!^~�v�5���|�if�5�*�r���~�6J������J�5rf�e�g;@X����eR�Rà7@���mG�8��=�Oy���r%&q	�����#\�$�,�W?�nXcⲸtLվ�9�l�od�S���f%@_1���@��{-n���-C�	[����`J��#�i@�F�8G�梙}�½����-i�r�g㍥�Av� Hn_�@�H3�-�@ԁ���Q(Է������~�i�nm+�@�͛�^R���yj��ׂH\�I9�8Rxz�R	xY]�ea
�**+mn���Zn�-����V���x����F?6b0����_����2q����9`����a�����Q��1���ޓ3�oj�j� ^��$�-�NRE6S3�O�4�b��=|ǫ��G�׻����2%��/�������]=�?έ��)�GGN;��9Ov1l�ﾝ^o��<�� ���T���@���������:��@Q���츘8���n}��1�ܣ=�a�x��T6S���k+� �ao�l�����<����.�ꇦ�0���_���菁�d��ߕG	��XΏ�|2{��/Bi���p߂J'6I9M:�m�̐��I b����z��W�R?Z�_ƌ�Ol�S�?da8�(��5��)�]c��d`8�ǚO*�N�ȉ�1V�W�\��_�[��F��wQa�}�f]���.�N񶢡+�.#WB�Ȩ���?�v���
c*��.��<!Q}}��չ���c���2�gY�r�IH`\�[S����;&��du̸>����]t���E��;0�C�<[�l��b��){���F�U�d#H8�s�Jd��
�"�D��y+�*!!��V����[��v��T���}�G.��&R�	E�,hS�vB\�Qơ�J��n��	ϧxZm��b�?�-i4���~y�w�d\<Na֠�b���`���Z��?8���?D�I�<�QG<a����z?��ƽ~���E2�P	�c����o�|"�e��#��8��ᨨ\{�C]�N���v5�����@��0�6���G��WV&i���}�!AC���3_�B�vHi�ٌ���!{Q�.��W���BA^8$	���,��\�CE� �2&�а�^Cym+����e�O����uv�,z��@bIR?��<�Mz��ELZ@DBbQ������u\J:�Z�l�A���u�	���ma����v�1����B��w@����X��jdâ`�̠�d��|o3�Ky'T���M�����]G�5��
����*�~�ga���ΰ��m+Ӗ��*��4l��	���~&#�pr��'���:�B&䒑5��$�56s�l}�PF��R�h��9%����
�֧��5����y.R垺8����u��zc��c" �Vr����ݬ%�EAr=НA�����ˁ���d�4�ݛ��g��^�׋x��{�q/a�׻�0F���d�8h/�^M%�n!Pm=������X(�_�1�̓��Tu�
��T/|ɠvR���/��7Qrt���,�Cu��R��q�$H�U���͙�.&-�9d�Fa˄/���!j���Ai�Q��tj��7��~����-1q����eK�?�D�h��[@�{F�ʡ�m�i��,V��!?]�<�3H�g7��]<���y�Z�c;�3�1e
EyF���FA4`���n�q�~�u�3^W�0!�q���瑆���$4g@�^���g��Ih^411�R���g��ÍI�j[��݃6]OI�:� <��#�}�6����~�*�X4�7͸g�m��J��V!h��� �~�2��c�J�&�� uI�|"ps�1ܿ�2��?�^�f�����PI�vĸLh�L3�y�m���N�]>�U�����ի[w^)줪Z��q�Xvj�gB�Hi^��!������I� ���q��"�t��;��(%5Cc+\���z6��86 �tMv��~��)!n��*	�q}|?��[m@$��E �ޡ���m_5�����}N�j��
c�����V{AA��湊�F��J
��!��r��o�9,8����V��VF<D)�J@Bi�zG!{��~{�q����Hl����q	��4�uU�8��w^~������@����r�'��.B����	v��b���_ȹ�鸁���R؆�ıޔ:�|���p��?fd��\��E/��Bc�����o�4��0���"F)�j	c���$�͂,�K�廸Id���S_��;F�$U=�⚚����Ӗ�G	��pm"��U��w}4�2Mؑ&�j��Ȳ���idb��1>�e��d���N�)i]�)mY�E�
޿��gQs�y�KK�K�|�A����<`NZW��E�6��=j����P����X��&)=�>\B�T&oiIw�*8��N)��`G��L���Л�ϑ�a"���XZo�:�������BkKX�G�~̆�������w7+���*�\┞�'EvJi�לk�S<��@�<q�OrT�K�'�9)�@��P��������f���43�ۢ[�n�I�͊��^�uھZ�
��?p�s^a�C���hJ,��}{	;���چu�5$�
]��3��V����0bKd����b{wy��n�|!��[��МV��b4= sl�u.M���I�n���vPB�B �g6O�K�(�r�
��Q�F��2�ֱYG��M��:e��ǥ�U��k��5��p�r��g��+ҝ�!��E�uk8}����w9n<�΄b FEE��_�M	5����r�c�X��1�>7�����&��3v����+̗��m���ؔ�e&]�����9�n��U
S�-Wޣ�`^��T����DuJ�)E�vy*��<���h)�iH[���*MM�`��H�Q���Y�sP�;
*q�,��?q�6|�z�R�21'RXt	(���{r�R�鍀@����4Q�,'`I��ߐ(F��9�y�Kc�C7G�9ۈ��G�j�t� ѐ��,X��'�QT���w�yr`΁�kn�	9��>I]�
�'���o�^�uS�A5��&X*���;���Yo�W��"N�����#B�79F�-��[��teP�K���t-�:�l�zx'���-�9��e��a��<�k}D�q�Q{@r0s����<��U��H_֝i�� @���O��ֺ�C 3��`;�A�1��U�W�kl2���]����U6�o�u+,9�R����)���Co���?B�+��o�����I��A���'� $1��Kx�.,%����)N2d�r��}���3�:�o2Σ����M����뻃�޴�=db"���"��1�� �w\TX�?� ��ݯuP�⼫DuvW\r2��B�����w���#��д��i)xO"-���M��)�i�.�t΁'�#w^�����wu���}sޝ�l�(N�B�S����|�x���Ͳ�0��|���5XBY�l����i�GY�Z��/���TwVGȁw�(cn�T�^S�kEp����&JGжݤ�eʍ�I���I<L(�;�S�k/�!� G�5N��F<xLZ�����ʅ��A�� �/������4a#'*�Z"�p4u����\�f_��
�ˎ�����F��4FW��ˊi<Z���ĺy�ڳ��������:����������U>)�!/;�q�4�����v�E�(���q�v�KaaO����v��g�\��soɮaw��~��gX��eXXh梻d�*������j�wB����+p~$��fG �\{�4._�ȪP�7g��f�����/ĮWt�9�黌&�+;!wK�~���#u	���4�WI˻��_����3k����j��D1��~��x�sk�Z�)��ĺ �H�L�[<oIX=���ȣ��8.�̤����w�Z��ïA�W�C�p�$�A�-����M䗘���w�����&&�M���?~$w��3�_=����y�=@���Ӟ*�),e�_�U�К��ί�Z���֊�n�����⿅��%�M�4GUZ�p�Tm}���˙����p�� \�Ez
���H�`�z���k��p
�?��,֍�cg��J0�@�ْ��� ��0��^*�^��bR����9���Dd�>����QL*蓿�0����j���c�D���v��a����?[q��^ε��'z�b<��{��;��OƄUv*@ly��Z5�.��X��al���tyӖ%Ї����	3�i�~-�[�c�nkۘ/�M�����O��,�q��y~���@�]����21aFJ�H�P�X,���r洛ߒ2��+�	6+��9K�Y#��_�j�h� �9.#��#�hn��T� .�-@у��cq�b��������c�v}W�Gp-���А@�\��d�'���DEi��=����.��b<
�(@f�C�0K��O-	�^�n��X_AJ��]c|N�,�979p8�r��aO�|�պ�q��0FQ�솭-P���~�%ר�<�"�)�`���۱E[eʕ[���3 �Z�e~�@Cc#P�@^�N>N@���P��;�-ѽ�st�#5b&�;�i�qD/�%�u�F&�r�5i���hrXJǞgD|�*��ׁb��x�`�u�
xᕌ@���[;h1����X�'B[_��������\`��/��Rn��\�oqu�>l�=�˩�0nys�������~�ID�ڟ(�lҟ���z��}��z}o�ʡzi7^���k�l!Q/n�A��S����M��x�ݒ�&)��Y"�׸��7Z��>����?�J�������L҂�����g�+ǧ��{�$k��fWr�[A�<��_`PP��e����q�9۲�A2�=#���Z|^B9Zn�;���D�P�AY����+6gH��	�/�.�s�~��*)�q�*����������е�����wp~!Y�3di��^���- K^-1�܈�++7�!��jD���P��r�������B ��lD�XX�4Z1�&̯E���,���
�r�vuDn����O���
�����^i�ɔ>D܃DXyz�~A=�J��G~�[`௪Ϋc4��e �9��K�KG� � �ԔR��F��"�Gݩ�셙/k�nmø	q�nkk���G��o��+l���0%	�V-鑾���\�r\*�2�?~Х�6�+I!{ ���Unq*��v\$��ќ�ތ��^+�Q����ƥ��'0 8�+^���������Q����j�!]��F�i^'��/���ӝ��D�ڥ�4gJl�@�[�nዽ~IT����Y@��@��/�0Ķ��ң����"ƶ����(ʵ@��' ɾ�\�mi �XV-_o��}}]��7\D��r�ܝ�⸪!u�z����`���a�]��Ԁ���;����9��#"B����2 �t��eYc� �k��+#v�HݭE�8��r�1�t����+#�؟���R�`v�h���1�ր�x0�뎫XR����fc-����:��XF�3�^'F]DN���顸�;3�֥�S��2Hj�T,�y��WS!�������"I�3^��#0p,�L ����_.q�V��� ��(�o�}�`W��`x���u�����|�N����@��7�\��_�Br��60��*���zxrg������
���8��@�|�ͯ~^۸#2(�����A��{k��f!m��o����	i���l'.�Eu"WFq���RO<�����OCdir�]�/̜���K��fT�H~[(+%S;�z����{�<X�>O����u�M2�T�{���L4�����HLT�|��)�ͦl���J����g��%<��y�꣼�� 7E���?�W�u���U3�,�%�T`TCs�~�Z�({�ў��[�7:<�}w�(����8A�Nl�8
:�}�1.�J������0����ea͎�.��#e�i<E�a���[��k�����ޯμѺ��mm�йl��V���f)��^������l�FX_T����;� �8��bwC��%^&n\{�M�x!k1�l*�]����3�H�I���թS���y!D�@�Df��|-�#Q�j���a����82ݬ��9tI�7�iy�@bh�%k _Pts 4O���|3.?h�]���u���R>X1���9h���p�UF�V��Ⱥ�z�U��������F�w���b������9�{6���տ���8�`W16�U�/9F`l&��}SF��&Ggp�����7�;�٘�=�|M�T7�r��l�ڞ$���ҧ���|�z�����)�2�`�!�vth�3���e�~��z�,(5�^�J6uƑ
���7]��Ge�����mr�Vm2'x�b?�NE��IHe�Lc;K�!k�ʹ�m������@o��W8+�I�*�i��Y��}�� c=�	��U�賠U|@�=b0&G�d��r�!�\��6�1kR�n���zH�':LWR>7���p�R��[��L�K" A*dS�b0���a���E�I&S�K�@��疖
���&�篖��vpjj��T�;��[��Hz�B��ֹ4��/M`�~�;�����E�,��#*��O���'�/�d��#����}X=�E�ѩ��P�u/N����50���fg�"$&n\��f��=��x12a����_k�xb<�W\���>�� 00Pc���> �f�����H���Sɫ�RC�t�g·v>9��`��_����R��½�#(5ՁJMV��� 'U[[{Nd-�Ϣ�����U��
��@�.����%aO33��͞Y�6�皏t!]ay����X�~(nط�G�M|�\��	��@�Q��ɪqwJD*6�+��XJ1,�8c�8����#^9S��ٳ;C@p�L�3�(B�P�!vw��)�A��D�Jn�k�D�V�S��9��̀�;��8��y���5�rE1�C��Ԏ��x{�-��[O���&k�]q�Wӊx���������������֛{� �U�J_�j����b7??I�Ü��p�R֘+��?�A��Ρu�"�~����4�Ab�`j�<7gͬ*8�ݨͼbHr�
͉.��F��ݩ!�D )ԫ��T4�d���d��r亰��'�Z8������K4�7 �}| Ï\��z�$5/����G=�n����I�� �qd2P`W܂�$1C�P�l�m�MJ���pr�f�+R�b���$��+O���2�=5R|�haS�Wa�!���XFo��XYd!���9v�4a��X-���d ��Yd�A�O\��+�������a(��N7 �!}Y�#��s�!�vb���o0�B��&S��7��<E�3���g��SP�J)E��?xX�1W��+(X�7+����L/��QZe�2W�c�뫈A �U� ��)�wς��:�2�	H��{�:cq��*�E�&��T!�ܧ�������K�YF��=�æ�n�@���ˋ�>��_�6��a�۬�T �����ZE�Vm�I�t�u7�'-m��Xu�	;�����7�iE:�Ę�v��/����r픭��2ņ�u���X5 Ս��\<٦��.�rEz�Miv����m7�{��]��'Q��9�/cs�t�P4S\r�W��`�<0RļS3�#�V��E�ǐ�+��kح�7���K������e�O���ÃW�b�0��[��$�R�+ԡ�#�eCn�LPh{;	�/��f��C��2��'{+q3�t� B�_�L���_�n��8��6$�舉"��T�ؽ�7��E]H�b��c��Xc"mh����k@�o��,pyޢ,��A��O��v����
������±��ح�
��Z�{A��.Շ�i�w��o����!�n=�
�8�>�ܿƍZW�(w��J�|�uw�w�u+��F�q�r�Lԛ���7�EÝb��y��	﵍5����� ��Mq��*A)		�:�ѭ�Z�^���*����ҴY�r5y�]�<M{m˅�K�0q������iKeڣpy*i6�ηR�fR�9
�݄<��MDEOC�1rb̖�_X
J�碧��/|.BO_����Ĝ,$L:�͌og9h6��
�ہ��Z1� |�j��|�㱿��T��1��C@,������ �_������;��'�6�o���g4�a�=�~��uCɸ�R��ed�>$0/��X)(��E`��lC#3��mx�K��D��N���E�'�)þo���c3�;�҆�a�^�|`&Z���$����0�[�B��x�uq�Ct?,:9?�vʢ�N/��9>��O�cNo��_=9�vj�����!�����N��=z��եo��c���A��_�z�1�a;��55��tP8r�3����|a���Y�wIe�넽x2j٢��Zrl֎��F�3b���^.��8k�n������E�j(��+���6�9Q���d:�K�Z��t�]��9�)R�]���l��hȁ�n\�&��ͅ��Nmj�:[��Q�so�\���q���8���N�wxk ��\�� 2�Md.��X���u5���=�B���`�5ْڊL�u���.�c�{��wP�`��3�����#�F����r~}�$�0�� �"*r���A����V��[=$Y���9Z�֋"��!²c��aLz,2�y����yM[���k{�Q��o)*{hR��Z�Z��+������)U��R#票(�*:s�g)�����ۀ�{s4�ڑ2�����׼7����a��盡2[u�p��p�4����f���spt�{#m\(&H\|"���Iql�XRZ#�L�ޤiF5@�"���̄�^1��L�3�>�4+d��2�;��3���N�pFw��dĮ�(6F��K5���X5rg�!{�M�d�ѝ)����r���O�Y�,<��˳&�I����$$�DBgH.S��p��I����	��+3�KY�$�O�b;'DT6�XĊ��T)��~z��1�GX�<c���^�9�`˶7)����R���M����b�(}t�g,��ԍ�~vΖ�YU���$a��1m��摟��,m�z/��q2�8H���}=X�~����W�ŝ���
����6��s��D�$�d�n5�phlw��	�0��']�G�]�t�C�!�J�$af�D�<�,��pYm��Wjܔ�������Ctp��')�l��� ��9�V���'C_�-�[t�-5|�V?e#=�5��㗥cI_�q[1
�=���}��o��(,���	r�ߖ,x3l/{kYm[C�䰨H����V�KP�hU+M~�J;u��#��7��7f���q��j
��2BҖ���TT���Ϥ������a��Z�G����j	o���;�}���h݈kƗ�{*�7�eS7�2��_ }�>QCh�淊��o6��b�\l�լe�ūq
��/�b��r=tG��Q��QЦ���.,J�ɳ���91f|�_4�c�9�pW����#$�K���V3{��T���Fe?���
��IU�h)&��ْ�I�pA��xl�ԫW�=l��$�0���R���W��lB��p�V�]'�%u�#Q���[q��5fҶ����v��N��cRҖe��}���o����}�	%��߸�<��L_p�بF{��B��e@��V�l5�z�����j6�zc�2f'x�"0�^D�P�d�?���xm��b�tay]�P��4�]�Uy,5���E�yp�&�S�'ڟ�n�#Ρ�3w]Uj�g_f3e�'<HOP)�H
�����?�@�C�΄���-����ی|�#���^�3m��á��'�Ʊ<�Qdu�n4T��iI��fL�&��K�N��>;xb~�#\<�tr�uuz�b_��H�q�F3;���&.���M۬�	_zh��cK�l�L�D��I�YKD?�p	�JL�^�SEf�����`fl�A������ܭU��E�b=4�-ǟq`i���X.�y655��l��Q!�Z��1������ۻ��5H�}M�Kڭ���=1�����F����Дv��4&D��0	v��b0�L��{#?vA�M����2�`}g5��<��� w���mU����x���ƭBI5{I�J0s,h�X��@����3۬|y���@��n�.,�h9.�\ׇ=��@��7�\h}�H;>o�jsQ-"HU-^9���M Sl����l��g��N�L���7��.))�T�$���K�cp[�.� `�!�֐���FU$��18���"���{�Y(Yy�N�W�ձ��=�H�7�a��* .l<	���I4�E}�f�x?3$\�.�_OR�:����,��Q��Ic�Hf�y����3"k|�Ԙ�X4�GpɍKZ��Q�Lt�9 ���V��+UƧ?��٤D#o�DE^�`�k���������D�T(���򼞿�Λ�:�В����1� @K�!�'AĢ���n�]Q�TG��V�-=κ9G0�1�ltV{��U��ts̝������r��O*j�1U���o�P3x��O�- ��� ���׷[��Qn��m�dc����"&����������z�'rK��ڸm���H���2w_��^���?Q��JG���m����|�$뒩6�/��̦����CS�oU[D.�V�w):�?��r�E�8*r_�D��a�י���Ȫ3��ą�6�$�����i�j�z�/O��&�/`�e�@.v���J�e���S��P�n�B�c*�3ry�L��2���u>y��[ڭ��{�֩��}ֶ}�$KP�-O���p(>�ߒ�ӭ�y`Fkf�����/%m��h���vpNz��o��3�j%�f��4�S�Ͱf dp�ٸw��,?V��+Nn�i���EeM�p$����x��w_�3�I:�cw�?!Ӟ����N�ȇ{~.c�ⱝ�C�2~.p���O���9;��?���'��m��d"�؊�!�-��B|gW<'���]����B�3�H��p��&���d3�M��O�k�-�8d��I_a��9���7h���!�pЛ��L� U�D�\��\����[w��y�b�@qq��α�Ds5MT6�𦜆/�^�_ #�za�Kaٕ�x�T��(���o�K/�T�D�A�߀�S�\0����eN����|�)�|���� �OrW	��.v��ĬO8]�@Da��R+\<�P}x�ǽZ�-M�[���V�{�d�Vͺ��&��C�u�f~�^�N> �˜u�S<iU`	���'`]�G�,Y�z-�@��+'�����Oӈ����)@��n��^�v��,��ٯ94`#ķ���1�2�Xu�F
>M.���$<�.!��3s wX��V��nd�������������KEo�Y�����b��
��n�{�"��>(��ׇJ�&1��0�ܹW	
���u��dW��ѫ#�`� s=+G�L�8 �f<"]:�yp�5+_~,��M�6Wi8>̧P�ɴ�� *�=���ϊ�	�cu������i3J�%-.��в�&3�C$��a��<�
�鶵���IYI�٦`��`X��F�]��S�:��Ǣ��-?�<��p�Eob����boQ������ƽ��*��[�i|�t��!J)T4wA��d�ǲ���;�bsɨBI�1�r���5t���h�O��c��z�����Q���T��	
�>����e|-�̻���$3�IJ�Ԙ��uj~����B�o2CӁ�f�h���5i*jD��4 F�%��%b$����c#�MHx(#����V�\x�� �+�Px���S��{�0d�-fZ�%L̇���Y�0i�r��#u��$��Ӆr������=��V?����AO���D~��)U�j�J�}��#��g�:�ʲd��������G*�y{���&����AG4������s>����
�/�eӊ*���t�:m���S��x7��lʠ�� 	�Ԛ�[��H�"ٍ7� �T1��t��K%���T���:�޿L��T��"�kP��\�\���Ш� �w�nԯ�?�"����� ]�W�FB)�$U�!$Mĭ��AY����-<g�d�ǖ���P5�sx�RYH3(F�h��ve��.ŝ�H3߫0XV������1�TU͞�d���Z�>6��*l,K��n5ׅ+_��3�.�r�����>0�����j/L��vI�,��� 99�*wc�<ω;��ۅƚ��l���`
�F�`v�\V�X#����΂9��Y����i
�p�;E��k�~Ad�?s�� h��>��.6��Y�){���?�qK��"٧�{xhaR�?e���B�����^n�8��߄�$�sW˔�}�͐��r����N/t322s�_�󲞵r�u���Wq�w�=�\I�_,c�6�<V���J����xt�/��°qʟC7�[w*O��uv���)��`�~���&�����iaI��=�V�pg�L����@zW.�UV�m/�9N��Vލ�y�C/q�����-;i��;;n����9������f��� I	�l��j����^��%�����ҕ<��r;��M��8��sP��9@��M�z��{�]rޑ"��&A8�m=m9@��
�hY�3B�����K^�%M@a�uy_�ዔ��D�����Z�Dr�6{y��BFs@Ѐ��D6�&VH[� ����@!�(DFnS�;󸢷� TՆ�,����m{b5��\8|�(���`�3D.�R01��Ah��!���<U�֢,qr�V]�ň�I��o �㐦�N:���3��+� F����D�1?�
$Ł�e����x�C����w�|��?������œhF@1�&g�����oW�L�_z�c]��uW�!�?��*	�M�U������W��B˷���l�ƭt�;*@�����#T�����۞�*��	���M���|����:/��K���r��:�]M1"b��K���D��$�g�F�m�|3t<�.�ԕ Ҍq�������GG.i�-���(�]y��V������NG�k��|2Z�B�]{_��(d��t��^Xn����(^�g�yL����r0W��T��G��<a��x�򢾆E��q����jY>���jN�*����M�F�f3z���'��Q����c)%V�=[���wN4��38����tN�uW������h~9Z��g�:ݰ�d������L4�g�kG�c1�)���-F�S�*�\�8������v�h5@���CKy!o��r0���M���39�vq��պK�񟿾$k�ٗ7���U�nˬѩ�>��u�P���w�dJ0���o��h`g�����l�������ŔT�a�m��˛�����ݼ�R��	�	��S-H2�'�;f�1YS�P7U@��i��Z�����=$���Y����P���p�Ѱ_�%g�,5�<��y���>޽jZZw��Gk��_� ��Ms������/�c��́�'u"=Ź����c4�3������A㟼Y˧Ȁ�ظ	��غ;b��HfS��oS#�_�h��8[LD���r]���Ό�2�9����S�.�	��������؄�������"���]�EҴ�fe���΀W� �00�q��>n�x0=��U���F��E3�N�T�\fDr�E�wX��؞|�1�գ����t��f��ݩ�;���t).7+H��#%5!R���J2��7
)�~�+�
����Qp|]O�Q2sotz��A�v�b��H4��y�`��:b��p�aV�1��1`�ӳ�M�"�� IG�c%�\s��� �k���P����ܹ�l�O�ؚD�.��t{ꠏ�����lE��Ibx���:�H8v�>��Ӌ��Y�D��")}-�5Gv>����d�Ѷ�8V��ώEO��N�w#kx^�,GXdv�[��Iw��6�􎳬|yݮ��_8�'����KUwh����dVD*�>�Qy:�S�d�� H�:]�R�~�p�����1 ��9�ne~�:bט�(���)�}܈wWҢM������CU��\��.ͯ�@�q����C%2�E��\0"�L���R~x��D.������}�C����W�x��Kn���a>Bn��}��bO�ўq�Ɂ�T���H������C���,�ΫiG�0�se&jtG�ԓ�M���~<>�hDJZ��'P���|��~I�Y������bt�jSp=��`dÌ�ǫ�>,v�<g_/��*�`t�v�p���^`k!��o2�w2M�����63���8qO�������6$�i�M�O���7�������i��P�N�*o@��RR����j�Ƃ/�2�C�b�%�ww���Y�����z^S��OB�l�]���aF�Y�fkك%�0��4̈���V�V' ��\T�h�I�����N�K$�z�=�/��gvK�-bf�,�b]��k*��`c+[���*\����l�n��]��,v��At� ���w̸��߫��yѶJ�6M�Tf�*6@_�$���g���}i�W��� 68�^�Z�c�63ԅ�7`.a�(���֬a�3^�_s�Pa�人�j-�S��޽��@)U�>��HN`�1�E�n���nu�wk�nN�{��*���@�>��ٹ\c�[4�z�z<�z;4S(�F��\���� (���WK�!�s�c��n��,�M +�9��I{�mT!���WJ�O�ѾI�gN�x:��R*8"4q�9�� �)�d�B�0���x�������߮(��o�\��Y�`n�$h�x��>�TOA��&�۵N�s�b5Z�&�M�ڍ^Ĭl�-� �!��ۻ"n�4sʀ����VB�)�l)�lx��מͰ%�)y�
gU�p${���V�����Wu��N�R&a�HY1߈�-~��ʴQ60�5��!8߈RiG�����2�ы�:J�[p�36���2]�zJ@��$�fS�<�QY>D4-M�.|�C�4x�'���'���a]�m��1���S��DD��K�{O��E�Srն�f���Q������Y{�$Y5hu���G�[@U�=o�G@A$D�AZ�n���F�;�SJPIi���n��C�p������{���\*�~gϞy�yfǾ�C���#ħ����T���6��;Z����) ��0�ʹ���m�B�i�;�I�N��Y�a1�~W�w��A4��p0��2n��
�a�X͢�P, ��`ӦD����iZD͓�-GHC�0��$�}Ry���� �b��N#�^s8;�d��B�<��,Z�v���=������x�P��9���@0��&v湣8�䌯_����E���QR���*��w�ϋ�@)�q�-O�	(@*��xE�{���+�� Qڈn�+?��`<��D�EηY'Y��ע,-a~$��)nA���!S���[]��C@O�����Ș{��Y��bO�Ҷq���jx���<�b�-3��S��PԸ��je�&'��fl[�?���>hN���o5�u��(R)�;��_�ø)n�G���H��	z�1�Z����ĺ�t��a�M�xf7g��еu�0U����mN@9���%z���W���
���	`��4a������Di����܇�0&���]���tG�I�Y�>e���(�_? ��"��o_�����˛u]�AԚU���gb�Y��_��,�NE3{v{��_Ț�����	/��e��w	k��z,N�kTRw~ZK�5���1�id�W�v�&N�l��R&���]/I���G0��N���o���3�}Q�ਕT2��9�ތ��!�X�t�d�^uމ��=F��!y���S붫�U��e�3�)��2_}�[�U��PT�	D��́�*�{����#폦<	
ȥ�3ߺ5�w��'���نe ��Ɏ����Q�����F�r�����ePO�r"AfF�޿�pks<��G��W�З]1�1KN�W�q}ʍm�ˤ���M��T���jAG4�g���:h�xz_ �
@&"��3'ׁ���Ggw c�V5�mk_,�T�4'��)�-��n�[�^K�����(!�B�q�|�Z�����fLu2Z��R����ͪ�:c;�VI4�����=�%�K���+q�%��E\���;��n��Lv.X�rf����=��\�b�k?p9$	����L����L&~��B�j���� W֘E�&���	�]�>�+������zz�o�_�^��CJ̏��:����$� ��S��D�I�P��|]����\�<�@4�%V.¦	V�@�W�C�vkյ�-tߌ��;�����e��&�p-Ԡ����-��S�~a��[F��x��q౯"�P@j5,�9�>�F*���+1���?�6��{�P�s�t�*��j/�����P�>�p�X]/m;��n�����C|�*��d��)�Y���L�0�="�#益>Kk���h��؇�� ��#�Ǥ��%�8+)��2�<���āz���$"j�Bv��aX�O8���?��+�Zh����ؑ�}��  o�]�K!^�$��X��<�rJ�(JeL�뻒��Nf�LS|LU�>8�#��:4��ļ�G��Ό��׳-	x{�X�ib�T���}p�qPu]��%����;�E$*iW��_Gɶ���(ҰI��¤?�D�/�:�S	��!�:�]a"Vn�v�JP�`A/�P0�x��h��X��N����AW[l��
Z�']��"LP�aH����uG(NT�`��pC�qg��k͌j�{��ش>t����hp䁙�ڢ����oW��N�Ks|�"St�G}��`���0���P�t�:�tE�W)FT����v:+����d��T�����w]���"{��a��WIL,>efY��_Sg����~��V^K����~�,�����H�ӭ��	\��Qg��f�
�_�9�A �Q N����㿠������g®?xѱ��HtG�|��$�w��r)�1�S��kIГTz�&������g���|�W@�ޫ3C��󛕐�_y��b�>��Az'�0��{z��hcQ���*Hp �	 �m7Pg�p?��9rM>~�@!I=`T�1�>J�;� xEL�CV��?�s�#.a �i�����!ꆷ�яد��O��XTq�����/\��5�/��ze�������YI�j�|(y9�G
t5�6�,���W����,��oX|���~r��Y�^�O8x|</%�v����`��q��ܕjW�1>�ƈ�ű1�r�%���|����1��D�jX��(�奤���E���ZܱZf�|P1A{����%�9O耨#.��BE�oy0:�tԙ�76�v5����c��A�	�����%���
+u�����	̽�Ř�9J��4�l���
��	������5���na#����_����@{��"�W��-��J��0�D���2"X����d�rz�:�u�8̒_���|Ǧ>z�t�u���994�D�L���AD�5�S(yP��W�F<]�j�b�7z�J1�yZ��B-ػ0"����*qP�}�#��-�5: �~�iQ�D�wV7��V�vO46�%X�LdSi��Ji��-��@a��3�������Wϩ�
�,��C��d �
��vlb͗鸝�j�+R��Iu��I�nc�UtQ�~�.�in��]����=w�����Џ��?�O(2f/��S��x���[����7a|(��L�+������߶ej�ϙ��P��� �>�'����W���'B�y#���b���M�s�1���d�oۇRZ��[ؠ5w��t��0�����|�G��/��gHO�]E�F�7�'%����N���Ӷ}�'9jS��/g}EV_��?��9j��Tx���J�{-�(�b�/Z�����u�|`�v�Q$2�ƷŚ7��(Z���.���B�_J����f��CD�r�͛4�G�\�S9)�{��s��QS���*G
@�!.L5���T�y���ǘ�j9��3�x8�$oxI�d� kSq�C|rYg��S��S�E�CA�"���G���GA�djoy�IW������?	��ۤ4�[S�%K*�A��D3�����~��Lq��%�������(���f�(��ʞ�b�v�V�n+\}��;��	���uU��{�#������+�b��V÷4��vD�`�c�]5]:�fgD���耭<�c|�Xwo�7WCB�
�Վ����x#����H�i�94�+�j>���P�H�B=F@|v�o�Y��".��
p�,/>��>��(,��BN�Gx��� C�H����V�g�&D-�Z�(��C�"E8�&������b������W}hC�HM���4��Ǡ� ���_m��ƴ�Q4k24⍱b��V���L�J�q�_??���]�J�"$�f�:F�V����T�m��d��Y�B��G��GC�<"�Е�K'~嫪����A�����~���\�����J��pkJG�%�  �)��~H�ƶӺJ�R'~ntRY��`�t';a�N�S���Z��X�����DG�[�h��@�A��IS�A>�u�+/�{��A��갴�VR��r�®#׫���&�r�/�������	�0�� <��}��#bJ�A���Tr��`�H�����k�ee�=cHxx�Q��(�G��}؍!��1ݳ��<�S([���j3vm���w����_H�~�&s��v�s��� �e*�Ji����h7:z�� �}��6�S�#1�$	��}��>��i��0@5czf��Hx�����:�~�������t��뽼�@/�V���r{�#��]���>���]M9Z���7���tQ`��.HẄ́J�N{�H)�i@�Q������Emഞ�֢!z�T6P�)X�;CņjH�|E�1�9�BL
��S�UR����[X�r���n����rO�+<�r�H�=�¨KWZ���Y�������V�����pF6X�&	6��<25vKЌ�'���Sܻ+o\6��QJ��6WP[�j�S4�S�d�n��,ˑ��jX�h����u��P�0ݣ�R����pQ�T���+@+��ГI���<at�`�((��nD
�}�5+U��?Sp����Νr�bF���v���W�%%�[��U��Ķ��q3#���{؍��!�o���k��R[����m��P��8&�i�ّ��w] Y0[�K��L"�t��B��i� 'eV��T��_���}�-9�@Yt����:tϟ��S?���74�	�0f�ϤHk���5B	����/N�v�y|����[+6�� �ͻ�� �Ff�\��邉���Ð���ÏPA.��3>rY��)�v�H0������.��!��k�5�N1�*4�>���p�D����Sye�k��o����oYW�b���F^ ���?�i�h�J/���ц^���)7���lx{��⍧A�mZ�?E���Kc���q0u�B�(��(���ۼ�nΓv��k몠ٟ�^c�;�����Gfv���*����,���u���U��,k[�GR��L��`=7����V�{��2���y���������/'<[�@�l�]ݹ/��fKFı����U�,�-�i�\��/V����$�NrTʵx%K���L�Q��óY���X7��p��&,�+V��T�U���1�OO�,�?]��� ����3�C���'���n
�7�_��U���:��%�؈��2d�]���Y��9��Ŀɠ#Z��v��o��B͟۷u�dI��!E(�}���.�%��$i���Ǻ�̿�&E�;�1����ű�j��j7�\�7��}�fH�4y��L���'ղ��?H��n�&�A�R��N�B��d�|��s����0o�Wwb5c�ݛ��.���[`\���Aj}���T�A����R���T�\�X���}�,q����#��a�`���DT��U�[�*��64dDߗ�ˤ��k�o��\����t�7*~+Q#��"$N��.T�U-����J�D�]P��EW啅>:������jO������{9�J�{�
��N��`��iN�F�[uu�]{)��%i��;)�̢�Ne�k�+�
KJ6q����M�
�p�/M� R5Tռ(�>�ű�O�E��5�o�u���«~��*�O��u\���u�?�^}�-�;�7_MwqM87r��.r�5[)BOi^*�74�����ԅ���6�1Ѿ�Տ^f���.�����R����{t������VD��m0���)�Tz3��ֆ����b]	$G�	�h����!ɖ����4��X�g"�8	:��c�د�G�/��;�$�=II�b�CP�"�=�L�5 ���A#ߗ\�85�B5^��A�İV�s��
U�^܂_�Y�!4�8����E�ڭ[��%Ϳ_:yH�%�loÔ��VO��H���bmlb���W�W����hn�[���ɟ�a��O�&a��bz���̵ͮ�l�'��CE��f���9��"�����5�3�lv�ɡ;FO���n�lU�����O�H���I��WgN�ކ�/v�1fe�3�aƶ轎�=���4�?��"�聉zm�)/�P"W7�d��Z�_���B>�qџ�$QEr��Q������-L�pJ�Ϣ��Z{GW=�~3�ٴ�~�����ԭ�>Gv(��E|���
�5������j��П��WQ�����͊载~s�&h;�L�y�U-�zY��m@�pMD�0H�	�\An�2�q4��V�~*�42��$�u�#�I ������ގp.4�=!�A	��O�uc����!����LN����H��� ��v�#iu~�6\<��Gtȯ��W�K�M�Ȅ,ǘ��{
t�6'8��&�/��������y���� 5��lи״���S�xúS�\Ѓ���qH��8�������>�Y
��ji1bL~ی2����U~�*�N��R����D���:�B��p))�Ž��^��&6�yAr ��$��'2�S��8��5ӏ�����1��]��cu��G�uj�� �O��'+(��(�ܴ\��R1�R�G�KX��q B�4�����h�$���8�e5K����0�q���T��ء���r���^�� ֋�&��tح��ᔅ[M��[Ī�ke ���c�.M�n1lN���;5�m������tRU�����F�|����Qi�dna���9�Q�������7��~k����K�c,+l|'�^O0�{5ԝs�\Ⱦ>�K_��x���ETP�p�8�bM�^s�888p;ݬ�^Ł��G�Z�S���~�/Q��6��Um=���$���b�gߣغ����E�:s$U:�ْ��*��R4k�5`���њ7���4��𑟐��R����&�ʈ����U�D���R"�����|�/�$T��:�#����1t���˨E�׹�' 
��P���>���3!f�j���ܮ!2L���l=b:j���̵�Rv��o�|n4��jH�2�I^h���3�����F���,x�\m>��ٴ�G��v�8G�uR�	����Q|���|���Mki�_K��NZ3Uύh��l�_�`�j��]sss{���4c2�+��̄>��`�'FCٺ5���9{��0�΍AQ_�>��n���r�Qo�9 |֛�?"�
g�a�0r��׆x�ծ!g*'<Z��y�js��q+�nx:|`}���h�w�G�>��,@(��T��:�Q�ql��]\~نf�0~-��#��s_{أ�����`��6����K_�g�����^�H��0{���2�4� �u�<7�N�q�6�����������2�58��v��B�OD���#tl��)�ʵ�_a��u۠��@�Y�ø�42���N�Pk�xZ8��ݫ�2��i� h��y��E�S����b�.��F��hz��ʻI5s^��/�M�6&����@8^
9����(�錾Pa�?���n�D��i���O��*�=�|=� =�袕(�؁�ccg�`��m�4$�Hsu�I�zO�[�=�j����R�. ��	� P�K H>��������V/���lR3��c��^N?��T�d�K*w�K�L8\ʝ����ǰ$!^Rg��M�uzK��`�����}�L�p���!�V?b��n�M|��&C�|�9�0���m�}�\z� R�����$�:�V@�l,/�m��݅ZI�q� �$#G�A<0�yMH�	��o��=5ݤH�Q���b�]�j;I��
��W6x
ݝ	Ώ�;�5ݭ�#�،/�%�>{�윺v��F	%?��(T��0���Ï���?V�C^���P��)��d�y )�C�%��E%�D��h()��)��j�S~g8�@�J�m��/���@�s;��z�߉�ϳ0s��l�g�ֵ+���j�{���!7��]~��|_����?���kP�S�-�~=�VQ�R1�6�	5m�5��((�:����T�����:U��yQ�s����'�y��n��}�d?Rb~�7Hf��q�uU$�L��lp�io�LR;����a#K����PƘ=>$7B�E�5��&�`ṑ�5t>��U��~.@w�w3�T���{���o��/�j.�5���9��,����w��������ﵷ����H�_�{C��{���K7v�ǖ�'(xo1_���"���w�&]x��S��"�2Ize��0�Z�,0���Z��WuW?�Q��.�e���Ы7��j���t�$;yw�Aw��"*X�w_�������ϻa��t�(�Qo�U�n���T����Kҕ�		{|�oV��:�L�H4�r�1�������1<FCs,�����h�~=zq����<L�NE
�t�tEݱl�^��w��ښsm�K���
O���	ը���(�xQ3BA�ﴛ�|�xڸ�[KY}b.Y������P� �{�'��Z~n�?�PY�@=}����i�a`�1p��Y161꒿�d�2�<���(mWFn?��ͷ�θ8�>h�wU�h�T��(�����_�٤fՊO�"���p�vM�w�wW{�L�M�F.ƩK:_xI�(ո#B�Iŵ>���D��#���6�|�ou�0�^*7��5�i�V2_��M$�ռ���8̈́��ۊ\����ii��Q@��R�"�����z�)�{���
���?Ek[G�/�]2����R�7lg,��.�jިI��[�����IJ�-o.̧��m>@!ީ.�X2���N���=�w)��y_�!/j�k,=zpi�̙�S�F�,)��螸�2�U�b2#��������Ӷ�ʯ�Z5��C��v�F��s^e�1���7qM6�'@��޾��R����n�\�S��"p7j;���QN�C�pq�N�=o�y6$_p~q���o�
���=&�D�y��N��o<������,e�=X�&�.U��K;es����w�n�Z��!�b}n+1����ר�7�#7@��In6 ?��A<����/�DF��6��)�K��~����S����(�^Û��R^�	xx3����ѫy�$Bc���?e�J�#M6��R蓤����O.�nQ���m#*��+��Q����F�{)�K}��I���"�3���_�XNv�aa1_�)����c4��-I<;���A���	�Ij"���>Y�\)���]H45��_�:�'���4�];H��`d��^�y!B$5s�i�����픲�w~o��H�38����K&���1��<�'�VkU���t��xM���)z�����J�܂Մ����4-䖦�z�ING0Ǚ?N��Д����4�`���q�H��V�t�zc��jr�T��q�6��1��!���β*�	^��k�6Q�3'�%K��4,L	|k|�΅_3�W��X�A�%�Ύ	&w
t��|����L)5T�Z��s�+�e��'�?)7n�ٯ���v&������E� �~�&z��}���|p��&< l��e�P(�zc����f#�-���_��È#�
�-"�*�Q�'1"пH�{��.����z��N�^�HC����QQ1?�~�8`v�O��,��s�����;T�s�	$9�-��:��Y�9�}�r�$%g�ޕH\P"���}�B����va��Jo�E�lӵ�vYX[���8���Z߹�9l"\N�@�IE�D-�[�~�`�k�c��,K镣��������S���������.3��IV.?b��X�^��MN��M:M��_!��T�?#�9���Ҽc3ÿo�M����ŶPy��j��3����u^M����G���|<*�\g S�dG�|�{#|y� �{H����)|r5cF̧k��1"=�#ⶸ{�_�(�>��^Pi�lU��y�]��MX�M�C�cz}�=�B�ږ*W!U�1w�]�������~�.�9ɧO���<�>����E��7��:�6����-��1FЧ�<)�3b�rY	�r�	�Аk\�7�������W]1��'}�#/5�輶���3���G�q�
�5�.sD��#o]�8��m�u��.v�ax�s� 5���.b�:E�)�e�z�K_,xw��{���'$�@�^�@H�֮��}x�Q��=���ӽl=�E<.�+���^�&�O�s�l���w7�ϣ��&��K�
��F	�I�[�LY������[/�v���cM�v1?�<�e�:w�Dn�tv�W�,ta�`ʏ�P�z��ng��Fc��%q��ߑ)6%�Ց�?���r+�S��;H��r��Ȥ��%1j�c���_�w�5E?��q~��i�oS}�����zc�FZ���G����p�a�6�@�C A�� ��l�����\E֌ݫ7�tȝNd�/�z��6�A�E!�򦢿�~=��|M=��ۻX��+��5�Xԣ��{�^�BܬQx�ܲ�.�廍�/
}������Ӄ=z�cwͪ�e���1�K���K6Φp���8-v�h��j�Z�i{�Pߺ���M���z�>`�l�U��kD����*�G�S�����p�|>l��e@:�NM�S���z��h�( u�6G������{�����s��f�f��2F�E\�>&z�i�Ӑ��}��������A�(\Q� W°�MA�^��U)�[(��k�*�U}��A�w��ub6�ޢ!=tNv2�����0:�Y�?5 G�"UG�&�s�(�;h"'v�OC�?����xW8�RLYLo�D��(f�U�|!O;ß"[]��(�<}vt:!}!��%C�d�:��jǰSau�}c�;�^x�vK>#��Z�?��4;����Cc���c���m_}�75�KQ`~,�]կ�6��_�wàOb��;��U4 �[������t�M�H�B�}�#	�tڣ��[*U��?�I#�EOЅ��0P�"�KRU�A�FB�s�c/��VY����nR�6��K2����~�"يHR��#]Ɇ��xsvQ
��ihƟ�O	��՘1�q�e�}Գ��n�mLP��u�ú �We/�xuƂ)��O��R��7����}M���H�В��_��bJ=5KKŕl��n��=�B��~Gr����G��+f��y�:�mj��X��y�'�:�<W���A�s8G/@�rJ�W11�F>�*˥��ջ���C/���31tvM��!@��!�S�!�<��',q��w�"Џ���4_���{ʨȸuڤ�Y��gT(�MaW��}#���xSb���T��Ź����ݩ���}��kT*��İ&��u���yZv���ln=�z����R�z���t�>T}��t}��(t��p��Q��}�u���F3�����W�����]��u���T�|�����PѝX?�:�zDz�+//�C/Ba�rs��0��XG���#�Ǫ�,'��?[���墖�t���l���ں�i6��e�ev>` ���#g�|��~5#�Nɫ�����D�%]O��������3�_�����!�Պ�V�����my����XA��ñ:�RxZ����8�v�u4*:N{�]j�b�Kg�������yI�^PZDR�z�f?�f���j�w�X�v��P\�\EAhBa�ؘ����v�z�����3�x,��A��;SILiQa4V^^zr������Z~r�f��wll�Y�4�r'���̵��!�҉���``G,I���C�㴁ao�qs�>��?��*���>?Et%9O���P�/so�5)J�gڟ�ijh�F�\x�S�'�d5Q���#��M�m6��D�Hʎ��b��'��+B�@��A�2{-.%%���C��f$���B���^.謖���>_�������5]����PV�����؂�}Ӹ$��F��_��Af�7f4��bN���.��B�NiLp˦��+E�p9����y]B���&���8 J
� 
'��{x=��<�bǌdG0ur8��=�������yƳ���G��r�7V��S
�Q�����o�F��NCIx������"��s��������9z}�<r���ȼ4����F]N�B'u$��n����i�/*�"�v����|7`�휬�g1r[5�R-��.�PqyɝA����l�|�}l�*$�e���zy�~��FNq��4~���Ѱ�q[��C�9db���6��/Ζ������k!�7�fT�~{������~�ݤ]ɓZ�P�>i�C���#�C�!�m�m��u�R��.�WY�k��2-��;�1L���J�y��˨���jĴ���z	CT-�A�b׌��V=bZ�CZ.��1��m�M�{��t�}�Ey�o��Q�
��n��A��t��4���9v5�ZLO�򈏋��Cc��A�%�;O�[�&�m:s���;��-����W��������9�H�`>8$�_��B����l#u�����˸П&l�+M<�A�'U4�������Zi����{��[7l���8/���m]d�>ݪ�_*Ot����h��&�s���j��r�{e���;hSY�OOj�F8�_R���d�H	�3N�uU�,�D���ݥ���*Y帄�(�_]o�@M�Ӗ�ԣ��E�����/�a��0���:^�K����S|��_���8	Ä�&i2'�k�jbJXz	��-����Qܦ���D�T���Ic�3K?B��oe``�֠��bNp�9Q�>nOճ���
����]]]k�O;�<O�N,��F��GW)CdF��sh[j������|�W]_��0c�΀��
�[S�l����LP��-C��Ⲣc��0i���eܦ��2�:�P�|�O��5>	�ۙi�}Q���h�Vȭ�#���7��0���!�/)a@�{jGq>26�Ѫ"߱��*�)aP���o�	�B_lwg�[��3�=<s͂��ۻ�<ք��+�+�pC�%�?�Q'��Y�C����T�_��hhN\+���r��w�~����r�)I�wb��) ����#G,�3@+8g�),��	� �>Va� 7L�Q���u5
�&�+@��ݒ�����Ƕ�u��`��Qضk�����#zT�'{���	K�)	ӹ���`�E��>��م��|u�QP��'�X�X�H4��뼊|?^��~KaT؇Ez[�^�U��;j�J�T"�c�����8�>���?i@>֊{J*�[]�5#lz0�&	PX*'T�	�"3i}y^G�b��ZC�a[�w���`\���g�[F13a�{v�j�N�t��V&w�gX�{O\@�P���k�pP���{At�?BC�.&��v����dx����+�;�nU�b�f%	�Ӣe�=&�@͛=� 
ZBO;B��\͸,·rMB�&K�ā��&v�@Z��[��Ɓ=�C���>܀�ސЗ���n>��}�톷FA,� �(��Q{+��IRE-Iag�H����m�-�sƭ:������}h[f˛ �`Mh�~m���e��~�"��5�~J�{���G�`CO��T��}(ݠ0ɩ.���W_��(a�O�y���t.�8� ��S�7� �00ȅ����	��Edx��Y����(�;:���U��T��_�*���*FT��>�9i]m�z�*J$��,{^"�:�!�/����8&,:�E��a�7����o�鶶�@�Y���tǣ�O^���9�ޘ�֩SF�l���B֭>�$*+#�@��.ݤ:H�D�� �'�hyݢ����By��|�a>��H�{�ë0�}�K���F�{��C�fȧ�PriĆ1Y��U�i(����,������Tm�K���}�|>�F2����Y���O��'lqYy9����D���Z���<

+����?({P`2��]�0&K�ǯL`o�����B�qJ�/zJ�?���)��D/�W�{�YC;|X,��4��G�!�|e�JUe��_Q1�m��Ey62���0�jvqC>+�h#�� n߁�-*��J����i
ܫ�kx���R�l���,Zo�3�|�-b�ik~�����5�)�F�G��#z�(��jB|��Q���֓ą�'D��_h�|�
��e�(((<�t��ݶE1Ѭ�bU������,#BA�S�N��E}��\�fw�&GK�D�gq���W����<������7pr�_�3z�L���<�B#���I
���l� (�I��S�.�iic8�}Ќw6f0!����<:[N����*���|k�m�rvu&��z��/ j���Q#�l�Q*��B��<u�ۗVo��=���n}���E�<�Ə����K���|Ÿi9^9��I��U�V����3�������k�~��U=<�S�6y���Py���bሿi+�n�f*�K�;Ǥh���Bjů��5peǅN�|�:���XO�E�Tg`�Mk��f !� D�ͮR4�EY�n���v\�Z��,��`'7�ɗ��CoT��	�@����׌��1�)4�������/�z��N�ɱ����0`�^�:�L]ZQ�ٔ0)E(rL f��r���IO��p�ĽMH��Ȝv]��&ޭ��^���D.3��Ԗ���\�}� lq�LF)l�K��A���<���1g�!��G��Ok���ƺ�?d��e�(d/T4�Zx���E�h�h�Ʀ�(5z�5ʟ6^�@���PŦ�_*��-�wA�b~8���R�z��9������ӿNЈLC��bSa��s�����'��X�>���Ǥf��+��O���fZaj��7Ԁ�5=�kn�?�:�Z�����������r�H�W�372(�^:9� n���Y�kUˉ����rB��)@��M����oOT]�̂�b��J�3����-ϺcP�\�&	 �ڼ�M!��9uN87���\=����HN�l�)�YdV�C�p����,��i�L��s;P���W�#�����W^7��Y�LfblLr���1�>MT��(���R�;₳a���[7w����e�G�hж6��kZx2���b},�we5��ʹ
6�N{նwD<�a4,�lכݐy�$�@���K+�Ö��Qѧ�D�~cSW�Ć��g4�����/]O9���YH�ǥ/��6�|Xh�%=� zJ~)�(j�4?�=�x�O�����.���4�u��7����n�&&HC[1�c5cv�-02�׺��{K3.A�`��w�5� ��  �
!��U���#h&
��E���vS��s�l��� $i�'�L�/#8w�0`��e�߹V0n�>"���7�O{b��~34�2�ck�fY68�&&�ş�U0�T���@7@�| �`y��Pa�~C* :={nC&��L�3�2x��N�鋾��<45��w�����.�!�e$yD�� Dx jB*k��8��M$j`��1�����qN��1?���]�mG߇)<|���tMK-�8_��?�6<�!��%��z��� gɠ�5�_�z"�#-�B3�=��.��EuK�`T���4����c4/������I�u�B�Cid���>W�N*�au"R�A�Вe��x�����Go���e$��e-/�F�{�1;�\�D�s>3�͏)�/�ម��{bgj��8��a���a����_����REJ��>��#%��xU���{C�l<��f{�� ��!4,ˍ���?���H?��5�h#|�aF�n)���2�gL�/�[P�k��SЊ��9� ń���Vg�շ%>�/�B��(���뇒���.E��"L�0N����/�����V�2Z��$����\�5i�΀T���$��z~^�g3���Ó�T5o����5Ѩm�%K=�DaݘOTv��|R�]�N[�������I�@T4������P��3z=�������,�z^�"}�녢v"ZX��E�̩�L�i����c[uA\@�E@9��7���-S�l< ��?�)� �Bl]��a�U8N��W럕�y:��dBəً��nVY|�¿� 6Հ�H�{BL�O&g12@r���Yw�h� q���B���%'��ÿ��l�;W���.)���Y���z���mQ8�w�L˗q0+$���� D A=���;W֡[�����g2*��
&�4����p��Wc`�*���0�����Lx�p��ˈ��J����;8�3tu���v��"Ns�}C_�[�Uq�.�a���5X�z#���V����c�(M�����]�S0�����iO�GJ�nKG@���a>�f�h���t	>ⳣ%�
xU��Ԗ�3,�����]2'9�-�K����'?������*jtA�v��1Ǥ-5�	�]����Z Q��ϟ�q��P�0Z]Ť��Yh���Y�%>
��%���5�0�=O����R�xw J���~��t�	���|��>�6�[넇��p�~�uVi�%��SR!zHV>S�c1|���3�K��5��K���f���������Z9��[�ӓ�Y?ߘ��E�F2��;��7����C�v"������+���kL��b"�P�R���U�,x`GT�%JlXy@"��oZ�_VK�;��a�(�+�ɒk�V������fA|r�x�ҵ4�����&twd@�W��,��M�����P���^.�Q8�����Q�=��1?�k0lF�M�T�n�
K.m��(��e��U]cҌv�7~݌���/��vǭ�&\`�K���\��;����J偳�X�8s��/-���%1B�i�M��`L��Զ�d3��B��B դR�x;�_��6�ͻ���2�ݽ�'�-\���@�b���L����/8e�S�����7��Fє\<�>�xB�Ь@�&P<��Dy>��Y�?�51F>`[Q &�:�Ʉ (P0�Mi��.�T��3}�qj4��evq�5�q�ί��Q=�����.�2B.k��>ŝޚ����P�܂��
pV���xw���3�8��Ye���G-��2z��<g�ue.���i�X��T��H>�>6_}H*^+��	A%2����~C��s��=>��uP���PdR1�ѳ�V�悋��$#%���Ia0�x�P�6;ȑ�Wh������s�(���;=��lGlM��ÖӽA�@/1�}(e{��ԗ��3���g��/��T�|nO���;�����q%ꕢacay���/#(�Iwo5Ir@)�˴�L����Lף��(�,}�PGn��ф��5�9*�O@~.X&�e�>Z�~B�U��~'��N8��(��`X�F��a�Cdf�y�!Z���5��XA���=VY?ӎ_p��[[������g�ךrz���V"�3:��_W::�cz�b%<vD�P�$�;r߱���G�)g���ڨ�dv[�)<4J��(����l�K���K���y����.(�535-��P�e~&�ۓf��wvV�i�W5���a��BXK�ZS�˞�d�|�>��Q=��7}�.�����Fy$��=�B!^�m;���iM��}��&�����n��G	��}Q`��mg����,*����ZQ����eK�Z�r{��)��7�����S�6�F꼉~�^���5A=�y�z9c����8�q��z~əsJT����db�1�e��3`wD#�l��u�m�Њ��.��CՈ/M�#""��DD�0Ê���q�^Y�uD�����-����Ub�#�p�<�k_�8o������o�\?x�ꪹt�qs-�!p�N��˂;� -�-t������~�/4��|�}�E%)X�<���fR��&��r���L,3H+�͙'��r�;75��ũ�\��Ϡ~� ��y��,)�塵�Ta��74��|����at��`��;�E|\�ܳ���+�2����| S��t|�s��}���-4�Pb?a�ps{�p�����0�A��!E�U��D�|흝���? �pݎ���+�ҫ��C��Lz�������gn��!��,s�:���5(0��M|��ɹ�]i�h1B�� U�A��j���=Z,--�)s���=��V�h?]��(��1�~J2-�^����B���/$E�	l�KА�%�@����I��4KJ�r<�=<��ͨ6��C)b5a��g�+U��{�J:��MP��dl��,6��bn�sE$��n�͵���)�R�A��%��XQ	����3*�%h��$I�E�A �	�"�Ȑ���" �� A$H��39	�Y��D	C� ��=z�{�Z���략�q�w�ꮪ�����̇)��yȲ��~Tz��/c��{���1f/��
�D�^$�^o)z����&�$߅�W���I�誮JӚ�|��Z�a'pS�FJ`+��~h����L�IظgŜH�pU�����~}�>�mo��U�|��uN���f�x�hڶF��mU��T	Hy��U�eu�O�Z���[��t3�b���o�˾��?U��]�8r�h�T��i�ɛ��2^��ct�6�q����h�63_+H��	8/栍��c��i�W���֜޽�E\RM��ޝ=:��ѥd1�:}�)�a8�3�����2v�����˚��.k�=d�)_����0z�I1�žX�[�|lqTa�o
n�%�E����7���x���.+x�l���Qp�;������QK���k���e�v��S���b��^��v_��{(�k��s��;��i�Y9��Jfs�����O�,���oŨD��1,`@�w�^�o����#�y�7	�ƣ���=�C�]z�����PCpK��A\j�ewuu|���c�����G m�g�'�$f0��Ǉ�S��C���3U�a*���X��;�;�|Q��|*�[�(M��ה��{����N��r�jiT��P\|��o�o���E@uav}��Qg��4��|pFR��N��Z/�z�L��p�}5G�b����
| 7��{Tn��݀Ath�<�l44Z��t��{�o�����#�ú��p�*H<�ͣ�#�x5��0�G�?���w8�
^�]����wym��G�{" _�kd�N��fE)8N�G� ���e/�!jv�<�/l{=��Q��px�(h�]�Q9C�B���`Vx�ڣ'1�
���������� Ĳ�pU���dY��{(�G��'|j�=L���- �a����*��wr'����I���&��9	%>�c����{D;ϋ��N��׈N���3���d8{�E~+� �,tZ�&Q���Z,չt��YP\�.�C�rnN8��x��sл�����G��
��⧲їN�b�~g��w��'�n�<:�kHezj,������[���:�Qosɗ�*0��MG�{������G�fmRk�
��	wa�+�������*k(���bޤ����'�@R��F����X�Y]�!�^jRj|�鮼���z��ư���y�3���v_"��@�6Auh1�g7�ѕ�qJ�i��.�>��l��#�G���[�5�&>75m�jvrT�$9K�#-�T����Ra+nM�5�7�r�\ᷨ ;KhF��Y_���P>�O.�7 ��O��+��S���jݯ�c5���Z/Yᚎ�'�:~'H��jQS�����z]r0u���S팄�г�������I�/'�'A�ģ[_�U�q�+�u�l=l��g���a�7��@��G�y&*r�D��f��%�6]�X4�Ո8�V��a���6�hw��33`[��A��|�d�.�����.� sg��t|ʿ6�w�'T�C�B�4�����	�L8>YO��H��q��`��κ�C\��⤂!�o�hL�،~N)#����|	�f�5��zY��A,�NԤ'T4>}��L��b{]�脣�%D������z����M^խ�/뮍?��-�K��g�}UU���sb_iu�X�֡)�3��ޕ��8BE���u�}s��_����%��k�_FƜ4$�7��%뫌���t���7Z}�ՅÄ��Y�'�	~K�gD��"�^���ۧ�rU_֫їe6]x�:L⇯5<*���qI��
S�>�a]
J�֩Q���%�c��"]y."
��W��\A�ձ��:��5�������_Gl]��9Y�A��"�G�
Z��_'yjv'o��]a��6�P�� ���:s��2z}BkD.����82Ӄ/�f}��/V(t�t�_p����782��$�G�So���앭�d��2�i`���2xĽ �W�=Ai��!�v�pɀ6	���[L��Ш q~ 4��;�S!���<�������������n�ɽq�%%����}�r宾�#Rb����ޚ��l��s�L�ѯ��!�_�N�ѧ�R;���hJHF���:����W5���H����yָ���� 6F�C�/˥�����q�k�h6ϊv� ~�իp
�_޻�����E�>�0��9D�[���b��a�T!L�~$Z�O[��^����g��j�R�<��Qi�� �J��h뱼��햪� ј���	�=+��
�������?�&���w�kц��:�-��[��A� ��>�4��w�RtT"z��{>N[a��kh�p�$��@g�`�ynA��ъ O
�m�
z	ϓ�:DU��'�?��dj��4|�� �sM��ż�C�H���4���tۙ�,����G�-��s:�K�b�5
�1g=�F�SPD��>�$3JQ?h&
�w^�@����D��i�t��k�U7�,F��26�.0��h' B�^�6Ho��M+�7����y�Q����po�O4��%$3֐�b�:{����e`�k�_@|�<�����9����L}�F�M��޷ۉ\u�-
v<�3~�D��sϾ\�B�c>mi'���u�BƁ؆*��X{�D+ ��;N��~�˲���bk��3|%W᱗�hb������v�
�J��J�)a�2#���iA:���0�3�$���Ӡ6�F��7��e�̕�W��%�����OŎJv��,�N)���^�8Ʃ��G���}PBٷ~�!��-�'^�/n�����τ.q���픇���#|W"B6R�l����("ū���о3���3��{O�o�llX��5�{�{]v�4�?�uh?�Ô�����yJ�(�~7<��u�+rw�f�]�"W������ m�3�B�CD��mV9�z���*1�����8�t0KPs�z������������$���h��_e��/Z���t&]�?��
/��A�=��H�d1`���2�������vy4�o��9x�>1_4�#s�[���!�bm��sBR,��@��(��
�����Y�֍��^Hn�����ce�t0�����
��[�y�ݰ��c�ޝ�Z��J���`��eR��5���ރ}�ˋ���a����'Z�qJ�|�/<�����m�|v��k����QH`4ʱr!/xh���%L:�6LN���YNߎ ���O��ҭC]	uM,\S2�\�v� h%s���(@���Y�v"���a7ΟY�@V���Z�O8@�)�s];��2>$iB̀��!����U����m�����^�����^�p���������R�rߟ�� jZ��:ID`���d�41��#������6]\x�a�@]�CD�
)�����s��&ш.�Kq��-A���	�x݁�
+9�H=�'�Z�<���Q����g�(R���cr!���]�JP�1X�D4�����iO�����+��7��6ל����^�����IQ}�Q�:ςōR{�O1%l��r��vx��;��9�~���cgm�Ѝ��SX��	m�|ߧ�����{����='�1�1=t,Jo�D�����~?��\o�>L+}aPL�ǂ��,�A�8���R���6�z���>��d��@e�9q���B�$��
G�Lߊ��$6�l�e��t�1ΖN�1M5��5v[6xK��܂���=!d#!#=���G�X8�J�~b���c�E[v�"�g����z7H���2)���4W�>F�xJN	�4���q7����c���3 ��m�"��(��JF�ӽ�C�_�H�&�oL@�0Q�W�� R�������hϱ� ח*�#�⧔�^ g�x7eI����3L]���Ɯ<늝3lA3f84
%�2���`���BK$"A���Ŗ=S(����ε�{��+��c7c�y��9�����L�GE��bZ�P(����#=R�2�y\��U��q�D�'[:>�`���Ď��|���z��P�k�>�E{Q�	5���VAH�t���Mbb�9!�,�g�x?��EZ#�`F��t�7{����� Y-���Ў	q@��h1zx�ݶ��T���� w_J�B|�a��7��4�~g��e`�ɴ�`<�9$������ý �|o~HBҕ��;�\Q�^ȢS=�!�4	[��T�X�6NJ�0O�{� �	�r�� �����+@W�et�RZ���a�l�K\�Pؖk�y1a����=�n��%e�S�5�?��������|@f��s���D8F���\�I�r�9s ��x�9���ۥ��%�<�U����ɇ�_|>MH�_s��B�>`��hZ�;��J��r{�L��PnD�8$j�'��R��]��ݷ7���@ʅ	�y��+ԻB�l-0�6�	w�p�0v�+�e��y ��Dq���Y�FN�6��7,����5�G�GcW�<���P8CG)����a�P=�/��V�๣c�}7���/�ޟW"�G���qUN�,@Z&����n�}�!G����Eց�i�of1L�am�Dv�_L�p17�z5�|,�?P�I��Ѝ�1�0WN�꜡�隘�|6��)=Wj�����
�R�O�r8yJ���zِ�<ZH��!WS�Q)����vJ�	�~J������y�I�qE�����7|�p�xˇ?i�E^N+�A���S�?|y^�be5�d�1��0rr=}h"���7�����f0x��a���9�R��� Pgc�.r�W&|��Q�P<À��%��"!ƾ����`,������\��qn�j<��U�;J�I��yK���27V灃�a6�#�+ ��Cy��D��������v�@^�d%�{���A�����q�A����YH�V�m7��A0���6�퇐}�!(��"�IP�o����z���fW��n��F�CFKN)�-<з�����Dxލ��vwu�h*bXz8����g��8���́_��j$��>�W�Xu��X�Y���$#�冝46�E�s�b]Gi7A��~�n���S��$�QmH_�}}q+&��y>Ua���@�q+����K ;@-��;�����q�pj@$��%��ݡ{�qP��,�*{�6�n����E+v)���h�ן��s�`bK�o�?���g���P�� ��sm��P�^83D#t�w�vi#1��~E�,�蔻���à�1 /�/�=HU#������*_(��*����|N�,���;��8 ��R���֩>Do6�5�^	ǈ��$bd�é⧁�������u�ش 3��9-��jr�#�y�$�.SC�������$a��I� R ���� �v��a�?Yc�l����x-jؒ�KBA�#]�$�#�ؖ�i� ��h�Jݨ��VL.|�Q���>��J��I���#��a#�U�x,�Tٔ���q~��n�#&���[ұ�V|�Π���0*��M#{į�����O����0�ѱ;S��X�����J�`�A��\DV��<��J��eo��Ҕ�j�ST@ i�Yn��V���wH�:/'���C��	k�����T�j&`TmQ�o� <ـ���¾�ys�HYǷ�%y���Bnݦ�W4v(�;�B�Z4m�a��A��8��s�"��\�x�����\#+.AS�Vq��w��+��W�5W�� ���t&庐bI�vn ƢTf}��7�y6������E�/E�kK̄IG����n�����oy��L�����
��R���g��+Lx��yU�9��0�T�8�0��LU��$ �$��5�CEZ�=#��ԏ�W�/����jAu"�{�_�n c�/n�Qa���dk~�H�1<����	_�ڝ��L����9���̛� �8<��͆\��qR�������u���>��(&�n�b8s����;��Ԭ��Q��s�Qs��2�T]���e����ϲp�N\,eT"t-�-���z����I#������ajsj�<
��Z��,�P�p|��<\R�����kK@,�Er�h1!]�'�@�(\^�>->���᧪������%�\I�����t��,���{wL+�֦�$�;~� 㹼�m�y�DLTx3���cQ� r���?��ҝ���o �_,M$��H�
�r�e,���-���`x��;�{?�	�ֵb�����4���Ο���}i�0���׋��dc����2�g���9��V�l��@V:}�q�>)H����1"�)��H�� �zUz�?I8�0݉�rª��3����yZB�� L����4R*�Q��

-ۻ���T���W5w�)g,�sP!`ԧ��8'����YV]���ԯ{t��% ��~]�+q�\�����@Anx��й��)��osPj�@F�4u���!�,� �w�����O/�p�e�2��-�,��W?�[��^sF������be��U��f�.��O��Xy8e�gXВ�bAA�Q��fC3��:S8�O���|u$v�'Jv(���k׸n�Z���`�Z86��ҧ;S?94XN���90"��e8�o����`T�������7��\B9\g����Λ]?�s^}����(G5/�I��9�_�枬�h�#��5<�z.���,��F���RK���C�<��H`J��K���$<c.d��2�@�'b6hs�0�ו�E%��n�U��n��R�j��
�$e'_��ǳ�Hڰ-�Z�jf�X�W�d��C�F5��NO��7��.��T��� ��>U��\<�|/j�"k�H5%���{�K@e FL��
<
�G�7bNTg�ϝ'�*f:��e��7�މ+��\�~�$�O*1�+E�4�Z�R���?,�:������H����$��U�������Ǝ**��ޱl � � -�m�^Vpn�c����^�ԧ���vg��ʦ��w�,6���)�f���5IT*|m��P����)�1���;uw?j��ŬhW*mg��5S*�8h��UalUK�ϸT�	�ΐ�����������ց�b����O��r�2#�I#2�Zj�Yc�vy�qlK� ��ԇu���m����YӃ��;�x@f��X0|f9�x��2m�  ;��5�Z��qׅS_}�\�r�j����j4��~{`e�܏a������_��.�:��꺯D]iH�A\�H=`e�+`r�1��_��P��甍�!��zUa@��>R�rsF�~�NFȺ�N���2��ř�R�;Ƿ��l�sk.B�Lj]x�B����7�n>jB�P�9<�0$��v/4�~S���L�'�m���ռU�r���aRT���;��Y��'�U���>��mƊ�|r���Id��Iy����w9����mEE��(��� {l�7�0�{#�K���6?�݃KEblN���(x���W&mh���a�rl뀅#.�N�Of����v��᛬�&��3���b�Ş��l��V�ψ+���d������b`@����m�7�H�����K(�Hr�f�0�ى�t>V).x�Ǚ�ҋ呆O4�!��$jFe5ŗv�.�Z�n*~����=,=j�� �=fx���V{&���e[�����iC��3�W`&ü���B���F �2K�KB}>Ƚq0I�F�y�)(^��#Y�:	�yr Q���k�d��u�*��S�jv!�u�tJ�Dd';��<o����d�4p�%fl��m���>�\Fakj��ۀ�_��5AO��&�ƥ@��,�O�Fp�qɷ3@�q�N>n'cr-ѻ�sw��]��cS�|�DzOx��1�#rLJxCd�ǉ*�
�|�^f��꜉0��`
 ��^�6S�6�~>7��9'(��x#l�;�gS��9�~��V��֝u�69m^������W�K�$��u{�45�XI����r�%��e�?BW��bs���G�`�^w-c�BP\$��J%=��ĵ0��%w�F�1G�8ȵ�A���E?8��-S�)Q��=�O��АĹ�3,`9.��t�`G�E�6�U7�A|:ՏB��:�+7-JC$�@��X�pk:)� =B��T�k��p��xH(8��Jب?�׼{@:��ܟ9���x�#�����$�ϱ-�a�Һ�J���bu�����3��|�pԧ���g���-�LE��X�Oy�@��8 ��=�9?�= ��<������Nv��x=���5��P�k[b��m��a��Ƽ-�סf⃾�Nb̯\����2<%�g�dIW>"��4y@π���������r�]ɞ=NiQHe������`�5dF��oQU�Bz�tՙkB&D���v7�跂U�G�;[�y�N�~ d_[�}A��(3��#�Վ���GR�G�D�a{��?�_[�� U��B�_C5����#/�_�n����u�ˉQY�)� ��A)9��?�Wb��͓�����Ub	D=�Ќ`7'*�n:~�5S�7�kPO�P�K+���zK�]��kCƛ���b47L�͞��
<4���x6�|vn���·����o1��VB;`��J�S8G�����ȹo��0H�
ei�^�P{z,���M���m��s�Sɂ/�;��?�f�'g�o/���z�����J�e�w8�i^���F�8���9Y�Y�[�����)m͘��=.x��&�p)<�NI�$�5rR���'�h��Wo ���*w�7ۘ�N�O��~�~��#2�~ܗ��U�.�����(J-����uPS�N�T�N���$O��M<}W@�<Ot�L�ą+,㷼�Rr����_�ݾ�0�9z������]�ӕ�y;��F�͌7)��C3֟���V���KOk�W߻3�1V�N��J�O���6'Y��6ğ歞�V�`�i�&��*__���� �!oDuVǒ����2���m��Ev��T���ۏ���'�﮾c���Z�2Z���û8��{��[��w���rhK�g��b|Y �[��K:��w�����&13>½y���M
!�hJ�
R[&�?m�v`�Y���;���n��JsJ�Ö/D�c�0�h������Q4�I'��Q���e'�e��^�Ș�t쏫uؚ
z�1���Wٙ9��^kK�K۪�~~M�����E3a��٦���E)$���r�'4���wx�_O�^�|i����"�����>�\ݑ�����Uۛ��ߖ�Z]���oW�����3���,��"��Ƨ�M��U���ӽ}�ӎ���cT�����ʳ�\��rP
���Y�֡�5��ġf��C���.���]��x:�Szm�K� ~+ʩlv>�zy~e���`����xK��1Mye�O(~q~,\:�⶛x�U��z�U���V��{���e&�qM~��{�ƾG��O�S;��ľ��R����;aʏ��=�����@����S~��f���7�3T�Wo�g�7��8����)/3(l��67�V�����<�ɷ�9��}�ϿH�/0�^�T�rqˍ����q���V߇�Ap8�͹
��?^����<3fr;f%|�B�E��2��x�����a&ɺ �� ���E�]'|q���&l���
q�Z�`�����Mݧ������>��Ӛ`i��V��A��J���k� ��͸~or(Y�1� �k�At=��Q<j>��Ry&"�9�2RW���_�������
;g^��>J�)�9�@��UEE���-�����_0���~"��<m4a�Д܆��la7����j]В�k�n����T�c�5�-'�x�sxҪ|u�9D���ZV�Zv����m;�A�>�3PD�0������������`�%_�U����7T���vX��G�M�Y��u��	P��o=w�!�A��[���v�gVsgS9���O�@�'�:t�ͧ�e��g�h�^��4n�;�3#�g�t�P��i
�XB,���-�kF��j�JA(	X����Ũ�KV��խ{@���{��N�F�R	!��@�!)�B�~���Ab\�i�|�������o:�yH���zMh;V`Y��
tL��
�=�K���MU�jw=q%�|��v{s�J-p��'� �;k,�S/��%w��P@��߿�xl~U�� ��%fI�n�~��E����S2��c�C�.&mZvK��y6�<:ϣ�� �/ ��{{]��˪M�3�Η������.�� _�|Y�� ����U��C+��!'���)�d҃@PmL.]�r:�Q���0�2JC7�ʶ�c4/o=h��'^T��O����۠Ո����_����Op	/-[��qTUъ�I�܆�P�}33��@ۛ����C!Wc��Y%��m�ZV�eݰ�Љ�Ƙ�T�"��d,��=��E쑊H��׮���c~Os��4�Ñ�� ��@�#~�G�F9�X_Y1
s]	�.��b�8�#J��c�W3%��l��?�^��9�<��H�9�ꂑ\B���\(�)�Iw񫃉�Y��s� t�<d�@�m�U�s�bZU�fj�q]�?��\
&��=�����A({R:��CJU��Á��5{����_��	_~�j�.`��i9�Å�d��'��g��'cN���p\1"h�Zo:�l?<a��f����M�U�Տ��l��bs8�4���ߊ�5,M����Ā�*u�����\�(M�����~��џ#(�l��h��8��d��f��K������rqjz!� 
���J�V���$5۲�?��X���U��III�!QSԏ�7m�5�~S��^s�r�߼��I�sk��f��\�n����'
%�S��Q.���[7�Alլ�������9�g�ɬ���_#�2x���{'���pz��Hn�S�B��Y|�e� Ŕi����:��k��7��� i޷Pg���|�|8�ǽe�a��	��G�6�t�m�����=pum-vǓ�����ÿ�vx����ۚ����6�_�J��.��$�w�=�8CE��8����8���	�N����3KQ�cw[+�A�Y���8H�������O����?�2U(���rCi�->2�g���� �VjE��'�n��H"sH-{&��E\�Q�(�5�}�ڱ�������YΆΨ������MM�0`��eh+�/���1hy |���%U��
���n���1��R#H���.�,𹴢?����dk�g`E��<�~�6�b��*|}*����5�����Z�0�EΓc�?�5]�o��A	�Ĺ50h+jRO
�'���\W��,;��Ȃ0w�����r[���z����!���݅�wC��cx�Q�W.n,����^�@tDè��ִ.vgx�^H��JYU�÷�<d���*���/㜹;v����c��@.��ے�%l�V	i���F"��q���I���t�XrtI�%�X���a�F�3��5���T�f=�4i�x��{R����_~z��?8H*m��O[M�O��-�ez��̝��vM}X�ܰi��|Th$��RI���	V���G� ���@נ:Ipik���i�����̊kO�L��D�rԑ-�T�2H3%f��ڿ�z0y�5�5{2Rb����v����N�N��K���7�'�� N^`�w4,t�$Q~G���0H2Rq+�+7�#��0�����-��xQ�`�IPj��1���[P�n��$��#��j:˂_G�b壝	��;K}�ݯ-����OH��S5�4V�b�g�/ki���T���(T�{��|��W*+~lϾ�@��p[��|����}r�;��$%�Q��(���V^�XC۝�]!����A�#{+Z�������I�kQ�Ѯȗ#uQA�r���R���@\��S�Q���o��3�"[��.DUe%��@�5���V�ZZ`�m�iud��ap���gGw��	�w�gnj�p���L�B�e�o,�<���=�&�RT���eWƈ�IAyL,4*�Y��e�s������K���Fn�j�`cY�Q���&�:_a�h�;^1�OY�9��2�V�K�[t���f]׳�d�|��W'h��)U�����x��Q]� 5n1�yG�{#9�ۣ�a��*��Y|��ˎ2�tq�g�d DJ�z�H������8�$�3��C?k��fyG�D�PVB�i��c1Apő�i���K?1�8�/�/m-���z��)��Eݛ�RE��yx�:�~�OE�'&�뤠�$@�h�Ղ��w�q%��xh<����c� �I��x�\7���dd�z�Ob�6�Q�b���v1���$j�q���PΟT&Պ`N���D��������I�i�]�xj�����!�I��(@�ki�߃k9�G�qR?�-��z�l�ݟ>�d0b+�����:�⺿Z�o"k�T 委�������ȕ�����(��I�F��1��QO���P@Ŵ,�~?��5�՝�|�y��2�ռiun�A�Қ��x�n'�_IQ+�54�!7E�R�xӾ��Epj��������Z�Xg#�׉�S��t�^���˿��� E��t<i,~��m���Xdnrv��J�-_2��9W*�U]�e"�G誓�-=L����G�]���Ð|�l���Z]��_�$F�b'd�@м��������)���KuS̛DM�j���^ײԞ���	�;�=SmuG�uA���_sT�֍��չ�?�6F�^-.6��d
I��s
����)O�B���L<*���8&����҂���*� ��~�����ǅJ�O�Vk�b��楚*� ��3 F�?�������^�[�H��W�Az1��3�H�n�%W��t�������p/
h	v�;	pR�0��'��ر|\h���#�ў�Wy��zhΊ���4�,ɶ'I�S�Ab� ��{葆�����=!�%x�y�̒ӣo���i\
`'ƕA�8�@0������'	�����2-닦�3��*��c��~t<B�h׆�`c�/U��!���=W�a�p�-"��E����W�4�1�M|�)�:����7���5B+;��6�JsT�V�[*A�!��Ჩ>��O�o5���:�Vg�H&�(�(�&t����8����)ZirW�>A��Ty��hw��5j(X������ �RCP(�ɫ�8s��(Zފ��LT�F2���Gc��^�*ˮۢ�$j�kh�P�-��JM��q��ɱ5(�w��)1�5�g
�T:����w{��r�����\r��a�"[�.K �����s}�MYY�W}b����CH����猒g��%�\V�����w �&i�f٭���,�	�R˗���B|1E0��W��/h�x���R�5w�fjc�x��k_�
d&2J�	Y4�G�Ԗ&]}^N)b\+�v�'�������x(b�x��;IT?+��BpJ�K�o�u�k�P�	Y��0�^��قЕ��k�����YC�s- ,P��{	��N��S�Ζ�6:�v�Ow�J� N�~ѕ����D���,ud/�Y����2�����2s���7�����	Vm ��t�ެ߬[��o��ˌ"e$�	�ʝ|.�]���?��?ҵI՞�\l؛� @���+H$2�h����;��P��� ���"@bm'��N�":�y���`�ر^��b�j�9��;�/��[ֺ,ݯq_��N���ܧ�e552nI0�w��7�S��ÇA^��B���7��f�qj:v�X)�jBE���O������KjQ�{L"F|~G�5�~�i�ai��d��s�T����=��u���b��FB pM���ǂ,����-(-;�h�w��Ej�������D�ɧƃ��U�x
�I�ˎ�4@S�[��":�'���8|���8՗y���I��v��[{���F�$�}ѥ�BPr���m7�YOvyo�Ɠ�0��	��?��a��Xp��T�P�zL�>v���g�ݾ u�l
%�Ǐ�ox�.��y����ɩx�o/r�Mdh�Ȉ��@*�X��-dR��聗t���ǻ	2�JZ%�����:N>]���J�!1~W_M*(Y�\R��e�Y�bCBsj3�sKS�[��	���»#�0�ǔGc��
&@b� L��t�H'�c�AQQ�4�!mIǭM
���@��ȟ&oXQ��*�ׇw�9�\�IQ�L/����$f	�ʝB.�]�#!�he��f��D��{���b��%/J�A���-i�5N6��"���q̈́�˟��ͺ&����9��Ĭ
ǾGq�ZRAз��mrh�!v#0��^�����g�����mxY�v�9���/dfĥ�#�5ʃ���Zثg!gx�B��P����E�jM��x�k�D|zX}�(a7����b�]��;s��	�H�L��~��븿�ZA�}/��Js��Xf��2k�d?���عvO��E��x���A�B��]�^�7x�!�U�����
���krۊs����0c���`�#S�u�d����<4��Lr�η�&A�*>TF>.j<����6�5���$\ ��g���XRo7��Ȇ���� +ؠE�uRn�M6�'9EL�(�7>�o9CaV�֙�� <�x��,k@&�@����[�B q�6�}�;U��j��8�����TR�4}�Ұ��©G��ݪ��M��aK�dR�	 ��0�#�6F��Y�Q�vcъ�6�<���|H&G�D�����_��'��k���y��Ȍ��`��<�'��[L��7i13R^ ��"f6�i��˳�Ch��#yڇ��spr��T8���qY�W�<)���iV��`��{m����|}�����;;�H�*��yS���L<m�Ƞ�m�7��޻�������=��V�i�Z${,�~���r��2cA{{mm�fѹ��..�SM~M��ǐA%#�_�~~M����kY����03����ktnC��0�X���-�^���C())	F����7��ć�&���D�?Cџ �1r2�`��1�7����$��o���!�L���L�of��G��J��ً�PK   Pn5[���7  	7  /   images/c1388d98-7bc3-4b7d-abaf-c89f09ba9dcb.png	7�ȉPNG

   IHDR   d   �   �\95   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  6�IDATx��}|\Օ�yoF3�Q�,��ލMs(� �$�e�%YbH$$�첛lv�K�Jv��@6� �$ƤPLq��1��*�eY��>�>�;�����k�Q!��~�ּv�=��{�}nFh^�����z9a�WU���CF8L�i��ϗ����;����ZI1�����r������P���w���|����N#nI�	�|��

���R��'(��YҼޜ^dD"T�����c����H��R����?|���"�����{?���ɳl���%Ɔ�g�� ^Ѓ��(���|�'� #�US#\n�		Ҙ��9�Ɉ�2<�4f��Y� a�WW�:~�}�~!�(��n�N�?@���p�SKR#c���q��!�L#5��������<�Yz���>�������~��a�i�.��կ|��:�}�gP8���Z��&�1�qAQo��:�bq*�����SvBOґ��M����6�8���Dx����������y��F���	G�=�ѼE����ڿ�Wzu]��B�r���ڞx� �P��X����7��{Ѿ��v����S����S���a�W 8sE��Hj���I$��O��1'&VP��	�Q]"q��*[�h�{MT��ǳ���*��E�u|�-�JOh�&�p���|���R:����S5H��'�L����#)����-4i3U�v;�1^|���¾���(�a�x::��>s��Y+h|�	����<��3ci&1A��s��1�z���@o0J5G��]��8�V���'WR݂	�9�XpX�Ĭ<�I3ǻӟw&:���i�o�Ty �ía?QwE5� n���;�8�?<gm�`6����x�=e��<��f�D輶6���'#b��=��$q�%��|�!X��*�y�8�����_��#1|߻�Χ�	妤&���`���5t��{��=@qJ��R���8��dP�������̪������ƶD1h׹3���)"a
�!�aW%㐟_��A���#���Z<�v�=]����q�_8ӕ�OO0�v�7����|�xJ��< l+�T1�c??Ε0���7��\?����'��ԆF&m�eDB������Y�ōh�ij���G�̗���d�� ��|��-|$���z���5�B��~���p���(콓�wx�X�<Y�w��z">&X���v������l�����1>��[�ƺ���Ŷj*�e�s��8�P�ڏ�n5�^nh��J��M��� ��F�->��D�{�4�tZ�cP{KW6�ԟ��m>���$�c��W���V̠I�mT�SW����U��B������$*�0.�~���7͝@�k�h|}k���DuǱ�Mc��6�	xw?a{��ml)ճ:���޾���Y�@M�c��I>>�W�����8���S!�W��Y/�&e�C8c���	��|��G��ڊ�����&�V�
tš"�T���-�*��_>�.���|,D��+��A�=�F�%���|�����^�:� '��c*�N�cS��l�	R*��q�1�X�l3�����+|��Q�}��I6��8:c��"L&��F�a
�M|Oѕ����զ6	�T� �cK�ag!ɾް0%څ� ��灿����ȕ���E��U����c�v0��ĭa��~������������� %=e~g���`Ά8Z������ =r�y�g�:�����y(̄�䷉\�n�+|4���a���+������N��]7D���� X��CA���<T����E7 u-�3�B}���)2�>X��8c�n�H�`_�R��~������rɓ�?����瓏i)�Q��'���\��;�=��}Y���q�S߲tݰ��w_B7-��o�Om���n�����`��e{�����q�:/�Y�ћt�B��-����nЧ�'\��fэ������!M��D��E���7�x	�˷���
>��~��)�o�����qVɋ��{�N�>V�����Yh��/a�L���|\C����'�Q�>�=/��"6�^�1�u���x�Do
�T���q� � >c�ک�+$Ɲ�>_G�X�'>���-k햸İ\Vx�m9=�vh%�G|�[|�Q������?��$�>$�!:��ʹ�K'�;�}�L�~�P�J2��':�B+�������o�6k�ˈ��������(D'�.qJHD�P{����4}����>y�L�<�L'g:Ts;5�LT�T �5��r.l�N�w|<Df����K�L㪼�GT���n��C��n=m�x�t����,�4Y�n�X
�?H� w�ӗ��SOp+�i1Qo �8�;�4��`��H�m=d������%D������*�
Aԋ���|���r^�v��N���AZ[����p��8%{Z����qͽ�L|�y���)��3���/���E�xp�$<i�?2�Vx���(�}�Ĺ�R�c�Î��N-mg��a�� ��|�W��!Nn/ ������
����k��8���bX�t�Ҋp9-�����;� ��QI]+��i���m��������y�#�}��z!f�����m����0P���/�'�>�!�Y�~SҔ}-���� 6<�����/��Ϻ�X��wT5���9�vQx���3T�R����·
.捗wr�ٟ�Z[��^Q7vd�0�ҙ��-��1�b��y��i��i
��?�p�;�)�:���0U1b�#2a���8쟶��*�Ť��u���#���/H�[Ld���B� �t�F�s��f�n�؁�Y~�]���G��)�m��ơ�+�w�t�3BZ�V���Y6��	���pt�G��������H{�d����@P�)����u|������w�u��W�9@Dt�{�H�^� _ ܏��Q�~H��z���V�(qS�����Ƙ���)���1~2�^��Hq#lrV�	%$�����<������J>�(�E� $j	���6Q/qS}��|��O��w31.��o��o�D�"�l0�J���Q�W��ňgq��$"5��;�S�<t�=�#�Z�����ȹ������ݍ�Nc� �$��8��Z/�Ũ`�b�|�1���Q��o!#�CU�.��im��	3���Yr��3����"]��c �2 ���MMt��3G<JUO>I������t<�>���=s���w$F�1�/����濕��Z��ߙ�Cp�j�i��w�{�\J��cL�	����x/��b�P�-_�Dw�d�M�L""�bǡS��&A�eD"},(0S�j��Fd"Ȋ������7Q�7�A�ɓ�\�������J0��L�o�C�`�i��)�ac*1ЇhԜ�@*���e��k7�!�Ik}���D�����H`\�z�j���9���I�g���������s����5�/�H��$,�ʫ�u�=�ho7��m��%"a�]�c�g�};�m	V7Ԉ�/���]'sF @�����Ӧ��C+��,�T/o�@ѝ�Q��������:�ٓf�� ߥ���x/��b�>�ڜ�P��Oi)�?q�~3ڍ�.F���;�N�.����Af }����(��ݻ��:��e.gk���]���������\��St�
��*ie���?&3��w7Sd�F�@zq�̫D�}�b��Qd�*���\��1^s� ;��+;x�bF����"!F��7)��0���2߇?���K�W_-�5X���=/���U#s��32�P�Cߧ�y��k_���]Tt�*������j����pO1sy�?��4$D�?|!�}V�Q��_�ĉRd���_����$�ϙgQd��>���P���~OE�>G��vQdӻ�:���Ȗ�� S)����
��I&z��vu��H+�����������C�E�=%�����~!����(�����/)v����X��T|�*���3kDJ=�S�nN2`��7	�%ZZ��	��?�Ǎ��믗� �����k)��� !�����s����3�S�&ϊ|�����"��Hp�V��Ѕ�s�i�15'Z)���;Vf��+W2�V	+b�U!
3g��&:;��ɧ���D�;��C�]|� 3,	C�����٭�,]JE�}�N^��|�]�}�O�-[��֭�Y���L�sd�W�B:sy��E���_�`;��ép���뿅 !�Xpq�=���	[�Hss����?�=����"9���3�a�џ(�Yx�����D��
�{V,��Dw���S����B��F�Y�D��^��xk+�� 3�a*��vrMO���L&L1+Li���r��l�э�^�o!ߕ�S7wXt���*�o:Jg,3;��EC��@���<����^��h��D8?��-s�F0h�%k����g0H���
Ah�+�p�v�5e��~´�軼�Ut�����1�5p<�Jl�~�`V e����������%!������L�ƪ�5e2^uK�3�g0e1K$@l2l3��BP��#�lh�qM� �T�p���g�Zc��%�׉�v����d=t:پ��/�H���M��n
<�8��kd �7�L1b� �w%���i�ݽ���r�3�.����0��9s��׿��~�-*��vv[�a��+�Z��8�[O�?��G��Q������I����S5Zt��~��٧>E�p�A$�A@D��?M�C�D-+�}���o���3�zR�%�BT�f;���_���,��$v�V���$8����k~-��
3���?�?S��=���̵��D4&��L�E,�w����\�&R�ݳOT!:�`	��T�M
1��}I�ld�&��X%D��g?�{`ü}�m�����>f�N���q�jk����pj��{�K��!*�=�?����X};�g���C�Z������a�B�>���2HE����C������|���D�Pi���Vu�-�0BBz~D$ְ��c�
z�)�����z����t�;Bk�&�y�����{�a >�{�)�|�Q�L='ׁ>��Ę5y�)e�^4ˣQ�d
 ��}�������ؙ��ѕ&�O�{��H�H{�m��5�\������x�lk,��a����ꚨ-���}�Y�}\W�C52s$�f�&��-�a	������_Hŵ�'�zƪA�'d����IC��3�`{�~��M�V�y
�~{�n����v? �h�w�f�_2�����	*
"!�@��|	zU Y��0�S���$�,GI nN@��Z���"uM3֕�+�$��Bq�v�&��牻���1!X��(x"�4�P��p��l���{���lOP��/�8�y���=�Vp�>gQ+�`6 ʺF�]�_eE�=�����S��C�ޟ��
?q5F��?b �����w�7�(N�<�}���Y�\p�WVH���?�Û9���sE5���Y"z�����b}�B}x�.����l���? O��\����YԔ�b�&��-���0��N��2�)� l�s�%�%aOd���zE9y?q���ih"��2V�g�5=�J�a���yx�!��	Q]ze�eW�d�e��{�=�B/�lzs6p�PG�B����F�܂eKMw�)���;�`]�[<��d��ʩ�oqd��. m�E3��bF�i���/�P�m�&������F8df��{IJ"pF6���lF:,�@�~�]u�E0�����d��9��k�¤Qrݖ�>Ÿŕ�>��#^*A�c�Ф���[���1�� �L��@�=q"�OQ��N�cNX���h�<��#��đ�L��O��z����X��#�n�4�a-����UO���A� ����H�W^N#�O����N���Ҧ�r�R�a�V`����^̣�.s��/Y �\�k�95)�YA_N�M�KЬ���%�(�̢b��.�WZ��}w��wZ`D*f��Xmt��C݋���4�c�V�Ӱ3B�;�	���Y�뚖�Q47"��̾s@�,��sG��^�٫R�C���3���'���:f����Eb�ٽ������V�u�����7�s�
;��X����N���X�NROd���(���#w,�p�9���zҬܿ����y�1�O%n7��b���6���,������y���7Ή �B��N��t��F&N�Q��?`H	q[����'����N��qA4ֿ����1�*5o���5���9^���t$L�m3� ��=̅K� ��$8Z��w}|�ʖ��� �7ꈼ�����o�����sd
��,RBD#+��m���*
��{�ET�P����z��ԩ���RGb��Χ�&�7����
����g��sΡ��J��'|����l�s��ℝlk�dK�*��e����h�Gd)A0Hm�f���:	��646DC5�Õ��R4�_g:D�kkIs��,O���@5e�:	@���M���BY�l*�7A0_�ѿ�$��F�ˠx�%�{�ԋ���z<�Ky�s�����Q\�� SigW��w�pj�n��F��|j�n�ڸ��q�	���--4� jt��y����jC>��o���K-ChNE�Yp���	:�͆h�pr
XC��wr �A�(anG<��~}a��6���A��A2�pc�k:�����hCv�O��gQY�NK('� �z2���t^%ܟI:���G��`K'$G�1�`�=�5F���!,��Ρ�g��H5��5kH?~�F���̧�˗'sjv�q�*������{�R��BFr����bAv�;`>�:�j+��e��<4(�NB���g2� �`�����;A��0����k먚�_�$�ܑ��4�6��@.���ʐ��:�{s�!���O�����q���	L���(����^�
G)4�F.o�|М9�cْ6Ĕ���#���F���ن�Y��9uB��{�+�RQ 0jwh���B�VW;�e�c�<8���~:YU�H���l�a#�\��O���!�A.}�%��.�K_f/��(3���,��.�褰cjD�1������j����J�D������:y��"�/:�*�a���Ym�Y'� ��A�~-��e��E�gL����g���X��4,�E�j�ҹ��y�2L��v�������ɱM�1,-�:&J&�x<�.��輣���O�h�نD#���!� ����fZ��ێ)j�~_�u�!lȔÇi%KA$Czc�C�"���8M<��8�&g�`<*U�	���MG�̦fr����8!������&M���ӓ������4�޸�t,eE �W;c��G�)9���,ٺ�|���Ce���U�s���3���߾���M��[C�-Y�u�jޮ=2��A�B�	���ul=I���T�);�Ш�!b�ZZh��Y%$�	!����5�M����G��Ժ:�8C�lC�6D
4j����z
fI�Ɔ ����>HA9=A ��kj�y�̅ ܓ����[�4 nj�8�6��˚y�`n������M��G�χd�h� ۓ��Ǐ��X۞%	�J)����L�+��� ���P�F]s�DI�S�Sg$;�N
����^C�z :Y��%*�y�|�PW���ce{��&G2�{O�SlmX�0�?3�eB?��nX�6�y���,zxj]�)������6�l�����OW�P.�}Õ���� �R�,/������֡ڃD�	����Vv���������zJ����(��@M5N�Bo�^�����ZH8[���gΤ��`'[�����b�AM�imU4Ik���,�.b��>q�"�&��`'��N�b�Z9�@͇�	�>
�8
�v��\��Wv��B�)*�Xl-��5����E(�Ӊ�2
g���sq��jC�O�Z��.���?������o�>;�O���5�J|b%<o���+������I�s`hھ��{�l�Ul=���1�Q*��Zl�;�겮�''�H:�{��&G�`��,vhtńI �A�DR@QJ@�y#Dz?��w�>+{���գ��z͊����+�<�t����Q�2��5my,|�{�b�7������pX��&�6e�; �����m>�Ae��_�6d4[/س��9Ҕ��ڬ��I:�� �#�Q�y�ԑV@�!�*\W|HM�6`���}�r��<O&��M��J���9�m�Y�����vT[Æ<�ti��^�*y�*��N~���j���F������4,c�B��-�^�Z�^Q�u'��(-�aY4>F�%����I�R��2�~Xv��|�_�6)���6dr�a��Jdh��]�tL}qȜ���ֶ{���֨8�W`�|r��/Kf�%,�P�����c��;C�{Zgw�;�a��>�6�v�ڳh!��L��u��2�*�G
0]�\�o�/�h<��Ӈ�|����*����{JJ�q��;�E�Ɋa��,+�#��l6$�ri�u^#u<Lq���Yˀ^
�e����Z}]�dX�cN�ui^�,d̉R��1������K9��T� ߊ�!�f�r�!V�u��o��b냳f��3ge(%5�BY�yK�������v/Z���:�e�,�>^]M{.�jC��*���"���m�渤M����N����:c����6D&ߘhC]q�l�s)i����[���G�e�N�{5*��GA\:M9�H+�f�C�
�N�e��Β�� P�}� �A-��)�f	�pGf����r�
ber���F,�z�+��6�����.
ѴQ��v��`�F��0�= �� ;�>��05m�7MN�&�����C^ÁB�����G�Σ��)V�W�����D�	�$Z\ZFnm4��/h�Eܯ�.r��V	�zZ��p�����+��#\36"*+l�,�����?b���#����8>��Q9�fH�qrw���ӻ�Dk>ӪRT��tU~�Z˨Y{����t`���#�0 �.��@�h���H	.ۋ��Z�H��ٔ^eI�m�z��އ%q��	wU��Ң;�y��?o��Pƹt�6j���]��}H�#-(*�g,�6t*���s 
ʒP�)<{�l-��2n��9Ѝ��8���q��N��4g��<��0��pQ@�bF,A|ظ��%�T�t��<�gj���l�._��7o���݆@\ u�@kiG�$���&�@���Y$͞%;0`Zy��ݲF>�4�,
�-�Pmb��y?��;�1V� Py(� Atkb���)�k?Azi�|�U���=��Z�H��CU8b�ԝ<g���ռ}�9�o�f!R����za�^UE�+�0?�mc|1;�k�ׯ����]F�>c1<F����N��j�L�|�5ʜ���+���R;צ����*��vM�DE7���Ҧ��.����d�d�	�FMo{;u}�:����܈L�O���Z��וц}�\C�R���l�w�� T�~�}�xy�=����������D��]`�u�7���)\'H0G�����:\>n�WϚ��|]7���v��7l�S{��n�*��@�Z�P������(�3]�()�(�8�i� ���߼e���B�4��*�(K�E�v����]T~�8Ռ#���C��< %DP�YJ��,0ԬZ����n��4�	�hJ���n���:�����tv�#G�K���ȍ�����k�MM�s� 1��'n:?�}H�;W���j�|������ ����tV���f����5cE�I(�>,*%��� �Tq`͞�lH[����ce�P#���1
��mjΥ�s�s0���$��VWG�`H8�8���b��YL��,|��Ã���.��j5����|�kٰ��|�QRF$R��`g��tKw@�D�j,�[g͢Mg,#g?��0s��C-V=,%+�=v����j���!*�2��T�d�� jj��;�	)+��j
��@��ϐƒ�`׸�K�P����{��7QL4�6��l����^�\UtC�Lp�=�FV3�8 �,Z�r7"�a�.;�q���2/f,���v����:����7n�;�E����Y���k8�"��������z1̆8}@<���fyY�7�C'NPp�:
bs�<|[^�Q|7�%huW%�b�)�P��[#i߾}t��!�:u*͜9Ӝ���ޒ����+)��z2�ج�=}:ŏ4�#�����5g���:I	�����.���E#���O�� �?]L@)�=���)�
����p΄P�:qlU��Y���)^W�j��q�d�y�Q��h�`9�LeI,�e�T�
�
�?�H;{��0� -�*�@ۭ��車EĻ2؋�n�Aqv�����>H����Y���^@KY�-ʷ�yP�&:uš�	h��O&�		���Ţd��&��˒�l�;�B�	7�o�e�"a��p�[����X�s����w���1�c���4f�'OR2���Q�w���O��Q><n&��s4Y�/wR�]�Ћk%���B[Cht��4o���{2���L�My���Y�S[G�q��2ॲ�-u"�̱5T~��x�I�iٝw����
����k�y�����/P�ג������\�,E�B�!�7��F>��Y��ּ�6�����MYg'Mm=��~v�O�Ρ��8�Y���U��R/&�ӟQ�%��;pPpe�Z?�����-���]q9���_��]K�^��B��#Lg�A��
����;�{�l|G���L��G��09�1�A�<��+�����{�Sσ�g�r*���Tt�����Te����Ý;Y�|����R�������k�3Jw`�>y�Q��!�EL�D��'�G.&���z�KJ ��C1�� ��B`�cg��s��;w����k���{)��0sri
F��쳨�c��~>S�ATX��7(�K$�}n���F�ٓf��
<��0:�M��Ә�-����T��������x�b���|�?����� ���|_L�W���l$p��暻X��{������_���)q�xaNy� �`c�xVQ���|��ꥸ���;%���i�JC4��#oi�8#����P�oB�#��~����{�:���i�y�����Tr�ߘ7YԿ�X{���S�3ϰ<��o��:o���iz�9�J��Vjۿ�쏓��>��>�Eo�W]I= !E�#8D�+�����処St�v
��2�,V�5k�w�%�3��,A�kx�D-{L:~$��Y�Z/�S���0��	�����fW������q财�]G�C����?P�.(��PF��1a�s��6m��G��� &���R�?r��_S��LXe4�<����Gޕ+����<I���}�~(��x]üf�?>(Nooo��ӭ9@�;E�w�Nzi	��Q��Ed�]�>L]���L�	��"��{^���4��ڿ�5�<8�zr�,����>�{!]#������Qb{����SՏg�|EX}!��Y���Ls�*u"/�W�,q�ȏd�Y�l*$��T U�� Tf_���@M	g+�P�>UqF.�:��\HDt;E�m2Ł���vpƴ}�y �рȟ���G@�Ӡ���(��L�F��`���e˖e|���:�����Պ�8w�9���U�v��G��=*jm{3 +'���}6%:����{	;G(r�4���1��( !�$���v� !@~ccc� ��ˁıcǞ��A�-�!V�q����DmbՂg'O���0##lB\�a��{�L�l��R�9<��N���/Ѩ���PU�OG�{�H:�*A2A���m;yk����Ǻ[�Dyv�-���.��^������ޜZB!�.��;?��+�Cq�BT6���
%!xǩ\X �ާ��X��Î�ʽF��6���{P���)�["33�@;nM�u���ܜ�ܗ�-^L��{� �5��QG�	�ΥJe���V砮�9県�L��YVVF�֭K8�m')S��>������s���ŋ(�E:��faI۱�%mP�N}���!}����)�d-`��E *�gb�l\
P��}v� �/�n�JBT��"�z6S�h��ۖ�`�<�e�Ξ��Y:!5l�&�-iÚ��K%Ghؗ����"�%ެS��`�Y��^�l����"H&.�K�N�BYBp�T��H
�g'����՞RY��)1�fV��2�,�dI[�����%��5ԮC`l���dX�,H�`3��t� qv	B]�N��)������C��x&]]�Ї�{(�u�ǹ�M%#�i]�\,.9� �q)@
\��3����T6�FM�"��_-g�{�祤���|N/@j�}���&��x}i�Br��ש��S�W���7�oFҥT�s)�+�(}o7�����`<U�J�����Ȣ!<6Mùt{���k=P�1�]v�,Ih[u�YN
M�n�7��"�l2ϥIɰI��RD��\�<*{`7�P7@�@R'vզ8_N��i�t��.��~�m��j�D��<�9Θ�jP\�ÞE:�*� �
�J�\9$6�|�;Թt�;�T�,�	Ik9��&k��5!z��a)%QHQ��>��RT�?@v���!�f'����	b�.�;�����U�ՕTM�NzY)�+�-�u�Þְ��sEEEI/Ǯ�q�~O���S%!��ȗ�@*��0bϞK�����S÷�"4�*C�� �� ��,��t{��)0U҉�T��7����.����ާN�J�����>����#E!^���`��e�s�:N��@d��AJJJ�m-����&}���̧;��#B�t	�'�  %!@��iT�0=S��&y
-���ZE��>ԗ"ac��Ϸ�j�tS'��v鱶?J�R{`�T�"�;�D�Օ�F���P���́��"����J���`�Y����Ц��t����L/�ϕs�	Pn�
L�m�b�\Ɠ��!��o�26[~,�34�Ȇ�Y�k֐�G���+���t	�E��v���@P��!h��f��^ַ�-O�K��������I[�,��wX6ȉ ��m�V��go�UT.�Xs�yI�B
� D)D���L�����T>L9 �7ǻ��S6v�%mu�t�ڬ�%m'S��!��9�L��͛��ߠ�3kNY4�S`(K�P�x�%mZ�%m
)�K�eS��9�.!��z&��D�@>2��6��N:�eI�o8�%m�@D*PϫWUʦ�l��ȸ�fP*��d��U� �d�*�v�fc��d`f��+P� ޣl�
���9sd������M�?��\jw��' ޑ�6�3��o .ׂ�?Gu�J�(ՔN�\@���V�Uvs&�Q*kI����k���c����}�*��VQeF����md�^�B
���c��� BN�8!R��(&��b�#S���իWӫ��*m�3��Ѭ�8f���^�{A:T��6-C`�0}�h?����s��c�F�5���Nr ��R ��<�N���3���U��Lv55�}+�N��+aP�ǳ�0_���n�ڥ�H��p^���}���nؓ���O(����K_,-�z��ݦ�H...����$_MMM2>���OGB *�S�9{�l��Qm�<�v":,��"�������J��ё�W����N���Y_.��
��r�����ӧ�;�Įfr���;A�A(`ҤI��ն����=���~��Y�b'�諲�\U���!@<�c�]/2 u�3�@�+R�J��ZDq�Hx,WuاWG�#�� ���qU�Ug�L    IEND�B`�PK   Pn5[�?E�  �     jsons/user_defined.json�W�n�6�C}i��M����)t�Ab����%bK^]6����$;v��v�ՓL���s�ЏA��v�YP.�j�ORg�a���E�������HQ���"8��q��^�k?^]0:@��O0����d�L�i��ԕ���IzS�Æk��:+�����Rd�Ha�Q�F�r����d�
�'�s7~��͹R�fT!s���QȔŊ�G���%&K�ERpMI"�#��rIK0����sO`�v�J߸?3�l˿���W�ͭ���$��>���ZM�b���l	��Db
�v�.���[8�Q� �\Wi�]�S{U���P�	Y��䟒%�DrDE�ɐ0EF!��������,���L/u���"x��N�����5���b��ϓ^|z �4���#����� n����^�O�|�N�{��~|��:v ��{�E?~T�C}�������E[�������x������x	*��Ou ?��C�:�z������Օ�@6�ѱ-f��]�T��c�q?AW�;�X�#qL�΀t5��@�H;���3tE��@�c���D?EW�{�=|����u��֬���	��l��2il��l��R�����:��v}�gev��5X6�>%i������}_�u~竴cڛ׎�b8�Җ��zɑq�k�x,;յcc)��!c8A<�ŒX�9!���aA6|�bň���Â�F���w�0�#�%aC%�HH�U�K�=X�x�����_��x~��e->%'�j ]u�>?�e��%|y2���;��g��g2�<I���+vђCQ�:\������U�k�q���6��ܨ�6���c��3-�ER$��=���[Ր7%Xo��S��צ�r��7B?�����z�Bm��*���0��Gi�I##��*�ʚx��7Z��[v��A�+ x��~��r��A�����+(�,�9�N2$�ך3�N`jS�jc,C�E1��I��\l�7���}��]4�h�w�:Oʇ����k�}�u�O��]B�]�� �~~�YX�,s7(���I�ۋ��-������F6Lu�K�%�0��d=�� �򯤼�xND�h/�u���M�U�����/��sڞ����y�)�N�:۝�p�7*���U����^ ���>��C���3��?4�95ͭuP�.B`[��c������PK   Pn5[I幯�  �;             ��    cirkitFile.jsonPK   Pn5[����7  �  /           ���  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   Pn5[԰�B� .4 /           ��<  images/44d6884f-a329-4b4e-966d-57539d09419f.pngPK   Pn5[���8  8  /           ��W. images/864a21b5-9f7a-49ef-8d10-822baf4f1419.pngPK   Pn5[�&�}[  y`  /           ���f images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   Pn5[����N �P /           ���� images/bcd2483e-cc41-4580-b81d-0411c3f5e061.pngPK   Pn5[���7  	7  /           ��$� images/c1388d98-7bc3-4b7d-abaf-c89f09ba9dcb.pngPK   Pn5[�?E�  �             �� jsons/user_defined.jsonPK      �  Y   